// ----------------------------------------------------------------------------
//
// Multi-Dataflow Composer tool - Platform Composer
// Multi-Dataflow Network module 
// Date: 2021/04/20 17:50:12
//
// ----------------------------------------------------------------------------
`timescale 1ns / 1ps
`include "../../fifo/fifo_interface.sv"


module top_8pixel_ms 
#(
	parameter DEPTH = 2,
	parameter FLUX = 2
)(

	// System Signal(s)	        
    input clk,
    input rst,
    
	// Input(s)
    write_interface.fifo write_port_in_port_0,
    write_interface.fifo write_port_in_port_1,
    write_interface.fifo write_port_in_port_2,
    write_interface.fifo write_port_in_port_3,
    write_interface.fifo write_port_in_port_4,
    write_interface.fifo write_port_in_port_5,
    write_interface.fifo write_port_in_port_6,
    write_interface.fifo write_port_in_port_7,
	
    write_interface.fifo write_port_h_alpha, 
	
    write_interface.fifo write_port_ext_size,
	
    write_interface.fifo write_port_v_alpha,
	
	// Output(s)
    write_interface.actor write_port_out_port_0,
    write_interface.actor write_port_out_port_1,
    write_interface.actor write_port_out_port_2,
    write_interface.actor write_port_out_port_3,
    write_interface.actor write_port_out_port_4,
    write_interface.actor write_port_out_port_5,
    write_interface.actor write_port_out_port_6,
    write_interface.actor write_port_out_port_7
	
	// Dynamic Parameter(s)
	
	
	// Monitoring
	
	// Configuration ID
		
);	

// internal signals
// ----------------------------------------------------------------------------

//INTERFACCE MODULI



    //DELAYS (x8)
    
        //delay_0
        read_interface #(8,FLUX) rd_delay_0_in_pel(clk);
        write_interface #(8,FLUX) wr_delay_0_out_pel(clk);
        
        //delay_1
        read_interface #(8,FLUX) rd_delay_1_in_pel(clk);
        write_interface #(8,FLUX) wr_delay_1_out_pel(clk);
        
        //delay_2
        read_interface #(8,FLUX) rd_delay_2_in_pel(clk);
        write_interface #(8,FLUX) wr_delay_2_out_pel(clk);
        
        //delay_3
        read_interface #(8,FLUX) rd_delay_3_in_pel(clk);
        write_interface #(8,FLUX) wr_delay_3_out_pel(clk);
        
        //delay_4
        read_interface #(8,FLUX) rd_delay_4_in_pel(clk);
        write_interface #(8,FLUX) wr_delay_4_out_pel(clk);
        
        //delay_5
        read_interface #(8,FLUX) rd_delay_5_in_pel(clk);
        write_interface #(8,FLUX) wr_delay_5_out_pel(clk);
        
        //delay_6
        read_interface #(8,FLUX) rd_delay_6_in_pel(clk);
        write_interface #(8,FLUX) wr_delay_6_out_pel(clk);
        
        //delay_7
        read_interface #(18,FLUX) rd_delay_7_in_pel(clk);
        write_interface #(18,FLUX) wr_delay_7_out_pel(clk);        
        
    //MUL_9 (x64)
    
//1�riga
    
        //mul_9_0
        read_interface #(7,FLUX) rd_mul_9_0_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_0_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_0_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_0_prod(clk);
        
        //mul_9_1
        read_interface #(7,FLUX) rd_mul_9_1_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_1_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_1_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_1_prod(clk);
        
        //mul_9_2
        read_interface #(7,FLUX) rd_mul_9_2_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_2_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_2_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_2_prod(clk);
                
        //mul_9_3
        read_interface #(7,FLUX) rd_mul_9_3_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_3_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_3_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_3_prod(clk);
        
        //mul_9_4
        read_interface #(7,FLUX) rd_mul_9_4_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_4_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_4_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_4_prod(clk);
        
        //mul_9_5
        read_interface #(7,FLUX) rd_mul_9_5_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_5_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_5_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_5_prod(clk);
        
        //mul_9_6
        read_interface #(7,FLUX) rd_mul_9_6_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_6_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_6_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_6_prod(clk);
                
        //mul_9_7
        read_interface #(7,FLUX) rd_mul_9_7_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_7_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_7_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_7_prod(clk);

//2�riga
    
        //mul_9_8
        read_interface #(7,FLUX) rd_mul_9_8_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_8_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_8_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_8_prod(clk);
        
        //mul_9_9
        read_interface #(7,FLUX) rd_mul_9_9_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_9_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_9_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_9_prod(clk);
        
        //mul_9_10
        read_interface #(7,FLUX) rd_mul_9_10_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_10_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_10_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_10_prod(clk);
                
        //mul_9_11
        read_interface #(7,FLUX) rd_mul_9_11_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_11_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_11_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_11_prod(clk);
        
        //mul_9_12
        read_interface #(7,FLUX) rd_mul_9_12_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_12_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_12_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_12_prod(clk);
        
        //mul_9_13
        read_interface #(7,FLUX) rd_mul_9_13_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_13_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_13_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_13_prod(clk);
        
        //mul_9_14
        read_interface #(7,FLUX) rd_mul_9_14_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_14_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_14_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_14_prod(clk);
                
        //mul_9_15
        read_interface #(7,FLUX) rd_mul_9_15_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_15_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_15_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_15_prod(clk);

//3�riga
    
        //mul_9_16
        read_interface #(7,FLUX) rd_mul_9_16_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_16_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_16_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_16_prod(clk);
        
        //mul_9_17
        read_interface #(7,FLUX) rd_mul_9_17_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_17_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_17_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_17_prod(clk);
        
        //mul_9_18
        read_interface #(7,FLUX) rd_mul_9_18_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_18_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_18_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_18_prod(clk);
                
        //mul_9_19
        read_interface #(7,FLUX) rd_mul_9_19_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_19_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_19_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_19_prod(clk);
        
        //mul_9_20
        read_interface #(7,FLUX) rd_mul_9_20_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_20_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_20_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_20_prod(clk);
        
        //mul_9_21
        read_interface #(7,FLUX) rd_mul_9_21_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_21_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_21_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_21_prod(clk);
        
        //mul_9_22
        read_interface #(7,FLUX) rd_mul_9_22_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_22_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_22_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_22_prod(clk);
                
        //mul_9_23
        read_interface #(7,FLUX) rd_mul_9_23_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_23_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_23_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_23_prod(clk);

//4�riga
    
        //mul_9_24
        read_interface #(7,FLUX) rd_mul_9_24_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_24_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_24_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_24_prod(clk);
        
        //mul_9_25
        read_interface #(7,FLUX) rd_mul_9_25_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_25_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_25_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_25_prod(clk);
        
        //mul_9_26
        read_interface #(7,FLUX) rd_mul_9_26_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_26_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_26_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_26_prod(clk);
                
        //mul_9_27
        read_interface #(7,FLUX) rd_mul_9_27_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_27_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_27_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_27_prod(clk);
        
        //mul_9_28
        read_interface #(7,FLUX) rd_mul_9_28_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_28_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_28_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_28_prod(clk);
        
        //mul_9_29
        read_interface #(7,FLUX) rd_mul_9_29_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_29_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_29_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_29_prod(clk);
        
        //mul_9_30
        read_interface #(7,FLUX) rd_mul_9_30_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_30_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_30_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_30_prod(clk);
                
        //mul_9_31
        read_interface #(7,FLUX) rd_mul_9_31_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_31_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_31_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_31_prod(clk);

//5�riga
    
        //mul_9_32
        read_interface #(7,FLUX) rd_mul_9_32_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_32_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_32_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_32_prod(clk);
        
        //mul_9_33
        read_interface #(7,FLUX) rd_mul_9_33_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_33_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_33_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_33_prod(clk);
        
        //mul_9_34
        read_interface #(7,FLUX) rd_mul_9_34_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_34_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_34_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_34_prod(clk);
                
        //mul_9_35
        read_interface #(7,FLUX) rd_mul_9_35_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_35_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_35_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_35_prod(clk);
        
        //mul_9_36
        read_interface #(7,FLUX) rd_mul_9_36_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_36_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_36_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_36_prod(clk);
        
        //mul_9_37
        read_interface #(7,FLUX) rd_mul_9_37_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_37_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_37_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_37_prod(clk);
        
        //mul_9_38
        read_interface #(7,FLUX) rd_mul_9_38_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_38_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_38_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_38_prod(clk);
                
        //mul_9_39
        read_interface #(7,FLUX) rd_mul_9_39_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_39_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_39_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_39_prod(clk);

//6�riga
    
        //mul_9_40
        read_interface #(7,FLUX) rd_mul_9_40_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_40_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_40_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_40_prod(clk);
        
        //mul_9_41
        read_interface #(7,FLUX) rd_mul_9_41_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_41_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_41_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_41_prod(clk);
        
        //mul_9_42
        read_interface #(7,FLUX) rd_mul_9_42_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_42_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_42_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_42_prod(clk);
                
        //mul_9_43
        read_interface #(7,FLUX) rd_mul_9_43_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_43_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_43_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_43_prod(clk);
        
        //mul_9_44
        read_interface #(7,FLUX) rd_mul_9_44_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_44_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_44_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_44_prod(clk);
        
        //mul_9_45
        read_interface #(7,FLUX) rd_mul_9_45_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_45_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_45_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_45_prod(clk);
        
        //mul_9_46
        read_interface #(7,FLUX) rd_mul_9_46_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_46_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_46_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_46_prod(clk);
                
        //mul_9_47
        read_interface #(7,FLUX) rd_mul_9_47_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_47_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_47_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_47_prod(clk);
        

//7�riga
    
        //mul_9_48
        read_interface #(7,FLUX) rd_mul_9_48_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_48_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_48_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_48_prod(clk);
        
        //mul_9_49
        read_interface #(7,FLUX) rd_mul_9_49_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_49_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_49_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_49_prod(clk);
        
        //mul_9_50
        read_interface #(7,FLUX) rd_mul_9_50_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_50_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_50_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_50_prod(clk);
                
        //mul_9_51
        read_interface #(7,FLUX) rd_mul_9_51_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_51_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_51_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_51_prod(clk);
        
        //mul_9_52
        read_interface #(7,FLUX) rd_mul_9_52_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_52_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_52_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_52_prod(clk);
        
        //mul_9_53
        read_interface #(7,FLUX) rd_mul_9_53_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_53_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_53_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_53_prod(clk);
        
        //mul_9_54
        read_interface #(7,FLUX) rd_mul_9_54_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_54_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_54_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_54_prod(clk);
                
        //mul_9_55
        read_interface #(7,FLUX) rd_mul_9_55_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_55_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_55_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_55_prod(clk);        


//8�riga
    
        //mul_9_56
        read_interface #(7,FLUX) rd_mul_9_56_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_56_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_56_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_56_prod(clk);
        
        //mul_9_57
        read_interface #(7,FLUX) rd_mul_9_57_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_57_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_57_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_57_prod(clk);
        
        //mul_9_58
        read_interface #(7,FLUX) rd_mul_9_58_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_58_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_58_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_58_prod(clk);
                
        //mul_9_59
        read_interface #(7,FLUX) rd_mul_9_59_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_59_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_59_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_59_prod(clk);
        
        //mul_9_60
        read_interface #(7,FLUX) rd_mul_9_60_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_60_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_60_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_60_prod(clk);
        
        //mul_9_61
        read_interface #(7,FLUX) rd_mul_9_61_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_61_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_61_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_61_prod(clk);
        
        //mul_9_62
        read_interface #(7,FLUX) rd_mul_9_62_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_62_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_62_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_62_prod(clk);
                
        //mul_9_63
        read_interface #(7,FLUX) rd_mul_9_63_ext_size(clk);
        read_interface #(8,FLUX) rd_mul_9_63_opA(clk);
        read_interface #(9,FLUX) rd_mul_9_63_opB(clk);
        write_interface #(18,FLUX) wr_mul_9_63_prod(clk);
        

    //ADD_18 (x56) 

//1� riga
    
        //add_18_0
        read_interface #(18,FLUX) rd_add_18_0_opA(clk);
        read_interface #(18,FLUX) rd_add_18_0_opB(clk);
        write_interface #(18,FLUX) wr_add_18_0_sum(clk);
        
        //add_18_1
        read_interface #(18,FLUX) rd_add_18_1_opA(clk);
        read_interface #(18,FLUX) rd_add_18_1_opB(clk);
        write_interface #(18,FLUX) wr_add_18_1_sum(clk);
        
        //add_18_2
        read_interface #(18,FLUX) rd_add_18_2_opA(clk);
        read_interface #(18,FLUX) rd_add_18_2_opB(clk);
        write_interface #(18,FLUX) wr_add_18_2_sum(clk);
        
        //add_18_3
        read_interface #(18,FLUX) rd_add_18_3_opA(clk);
        read_interface #(18,FLUX) rd_add_18_3_opB(clk);
        write_interface #(18,FLUX) wr_add_18_3_sum(clk);
        
        //add_18_4
        read_interface #(18,FLUX) rd_add_18_4_opA(clk);
        read_interface #(18,FLUX) rd_add_18_4_opB(clk);
        write_interface #(18,FLUX) wr_add_18_4_sum(clk);
        
        //add_18_5
        read_interface #(18,FLUX) rd_add_18_5_opA(clk);
        read_interface #(18,FLUX) rd_add_18_5_opB(clk);
        write_interface #(18,FLUX) wr_add_18_5_sum(clk);

        //add_18_6
        read_interface #(18,FLUX) rd_add_18_6_opA(clk);
        read_interface #(18,FLUX) rd_add_18_6_opB(clk);
        write_interface #(18,FLUX) wr_add_18_6_sum(clk);        

//2� riga
    
        //add_18_7
        read_interface #(18,FLUX) rd_add_18_7_opA(clk);
        read_interface #(18,FLUX) rd_add_18_7_opB(clk);
        write_interface #(18,FLUX) wr_add_18_7_sum(clk);
        
        //add_18_8
        read_interface #(18,FLUX) rd_add_18_8_opA(clk);
        read_interface #(18,FLUX) rd_add_18_8_opB(clk);
        write_interface #(18,FLUX) wr_add_18_8_sum(clk);
        
        //add_18_9
        read_interface #(18,FLUX) rd_add_18_9_opA(clk);
        read_interface #(18,FLUX) rd_add_18_9_opB(clk);
        write_interface #(18,FLUX) wr_add_18_9_sum(clk);
        
        //add_18_10
        read_interface #(18,FLUX) rd_add_18_10_opA(clk);
        read_interface #(18,FLUX) rd_add_18_10_opB(clk);
        write_interface #(18,FLUX) wr_add_18_10_sum(clk);
        
        //add_18_11
        read_interface #(18,FLUX) rd_add_18_11_opA(clk);
        read_interface #(18,FLUX) rd_add_18_11_opB(clk);
        write_interface #(18,FLUX) wr_add_18_11_sum(clk);
        
        //add_18_12
        read_interface #(18,FLUX) rd_add_18_12_opA(clk);
        read_interface #(18,FLUX) rd_add_18_12_opB(clk);
        write_interface #(18,FLUX) wr_add_18_12_sum(clk);

        //add_18_13
        read_interface #(18,FLUX) rd_add_18_13_opA(clk);
        read_interface #(18,FLUX) rd_add_18_13_opB(clk);
        write_interface #(18,FLUX) wr_add_18_13_sum(clk);
        
//3� riga
    
        //add_18_14
        read_interface #(18,FLUX) rd_add_18_14_opA(clk);
        read_interface #(18,FLUX) rd_add_18_14_opB(clk);
        write_interface #(18,FLUX) wr_add_18_14_sum(clk);
        
        //add_18_15
        read_interface #(18,FLUX) rd_add_18_15_opA(clk);
        read_interface #(18,FLUX) rd_add_18_15_opB(clk);
        write_interface #(18,FLUX) wr_add_18_15_sum(clk);
        
        //add_18_16
        read_interface #(18,FLUX) rd_add_18_16_opA(clk);
        read_interface #(18,FLUX) rd_add_18_16_opB(clk);
        write_interface #(18,FLUX) wr_add_18_16_sum(clk);
        
        //add_18_17
        read_interface #(18,FLUX) rd_add_18_17_opA(clk);
        read_interface #(18,FLUX) rd_add_18_17_opB(clk);
        write_interface #(18,FLUX) wr_add_18_17_sum(clk);
        
        //add_18_18
        read_interface #(18,FLUX) rd_add_18_18_opA(clk);
        read_interface #(18,FLUX) rd_add_18_18_opB(clk);
        write_interface #(18,FLUX) wr_add_18_18_sum(clk);
        
        //add_18_19
        read_interface #(18,FLUX) rd_add_18_19_opA(clk);
        read_interface #(18,FLUX) rd_add_18_19_opB(clk);
        write_interface #(18,FLUX) wr_add_18_19_sum(clk);

        //add_18_20
        read_interface #(18,FLUX) rd_add_18_20_opA(clk);
        read_interface #(18,FLUX) rd_add_18_20_opB(clk);
        write_interface #(18,FLUX) wr_add_18_20_sum(clk);                 
        
//4� riga
    
        //add_18_21
        read_interface #(18,FLUX) rd_add_18_21_opA(clk);
        read_interface #(18,FLUX) rd_add_18_21_opB(clk);
        write_interface #(18,FLUX) wr_add_18_21_sum(clk);
        
        //add_18_22
        read_interface #(18,FLUX) rd_add_18_22_opA(clk);
        read_interface #(18,FLUX) rd_add_18_22_opB(clk);
        write_interface #(18,FLUX) wr_add_18_22_sum(clk);
        
        //add_18_23
        read_interface #(18,FLUX) rd_add_18_23_opA(clk);
        read_interface #(18,FLUX) rd_add_18_23_opB(clk);
        write_interface #(18,FLUX) wr_add_18_23_sum(clk);
        
        //add_18_24
        read_interface #(18,FLUX) rd_add_18_24_opA(clk);
        read_interface #(18,FLUX) rd_add_18_24_opB(clk);
        write_interface #(18,FLUX) wr_add_18_24_sum(clk);
        
        //add_18_25
        read_interface #(18,FLUX) rd_add_18_25_opA(clk);
        read_interface #(18,FLUX) rd_add_18_25_opB(clk);
        write_interface #(18,FLUX) wr_add_18_25_sum(clk);
        
        //add_18_26
        read_interface #(18,FLUX) rd_add_18_26_opA(clk);
        read_interface #(18,FLUX) rd_add_18_26_opB(clk);
        write_interface #(18,FLUX) wr_add_18_26_sum(clk);

        //add_18_27
        read_interface #(18,FLUX) rd_add_18_27_opA(clk);
        read_interface #(18,FLUX) rd_add_18_27_opB(clk);
        write_interface #(18,FLUX) wr_add_18_27_sum(clk); 
        
//5� riga               

        //add_18_28
        read_interface #(18,FLUX) rd_add_18_28_opA(clk);
        read_interface #(18,FLUX) rd_add_18_28_opB(clk);
        write_interface #(18,FLUX) wr_add_18_28_sum(clk);
        
        //add_18_29
        read_interface #(18,FLUX) rd_add_18_29_opA(clk);
        read_interface #(18,FLUX) rd_add_18_29_opB(clk);
        write_interface #(18,FLUX) wr_add_18_29_sum(clk);
        
        //add_18_30
        read_interface #(18,FLUX) rd_add_18_30_opA(clk);
        read_interface #(18,FLUX) rd_add_18_30_opB(clk);
        write_interface #(18,FLUX) wr_add_18_30_sum(clk);
        
        //add_18_31
        read_interface #(18,FLUX) rd_add_18_31_opA(clk);
        read_interface #(18,FLUX) rd_add_18_31_opB(clk);
        write_interface #(18,FLUX) wr_add_18_31_sum(clk);
        
        //add_18_32
        read_interface #(18,FLUX) rd_add_18_32_opA(clk);
        read_interface #(18,FLUX) rd_add_18_32_opB(clk);
        write_interface #(18,FLUX) wr_add_18_32_sum(clk);
        
        //add_18_33
        read_interface #(18,FLUX) rd_add_18_33_opA(clk);
        read_interface #(18,FLUX) rd_add_18_33_opB(clk);
        write_interface #(18,FLUX) wr_add_18_33_sum(clk);

        //add_18_34
        read_interface #(18,FLUX) rd_add_18_34_opA(clk);
        read_interface #(18,FLUX) rd_add_18_34_opB(clk);
        write_interface #(18,FLUX) wr_add_18_34_sum(clk);

//6� riga               

        //add_18_35
        read_interface #(18,FLUX) rd_add_18_35_opA(clk);
        read_interface #(18,FLUX) rd_add_18_35_opB(clk);
        write_interface #(18,FLUX) wr_add_18_35_sum(clk);
        
        //add_18_36
        read_interface #(18,FLUX) rd_add_18_36_opA(clk);
        read_interface #(18,FLUX) rd_add_18_36_opB(clk);
        write_interface #(18,FLUX) wr_add_18_36_sum(clk);
        
        //add_18_37
        read_interface #(18,FLUX) rd_add_18_37_opA(clk);
        read_interface #(18,FLUX) rd_add_18_37_opB(clk);
        write_interface #(18,FLUX) wr_add_18_37_sum(clk);
        
        //add_18_38
        read_interface #(18,FLUX) rd_add_18_38_opA(clk);
        read_interface #(18,FLUX) rd_add_18_38_opB(clk);
        write_interface #(18,FLUX) wr_add_18_38_sum(clk);
        
        //add_18_39
        read_interface #(18,FLUX) rd_add_18_39_opA(clk);
        read_interface #(18,FLUX) rd_add_18_39_opB(clk);
        write_interface #(18,FLUX) wr_add_18_39_sum(clk);
        
        //add_18_40
        read_interface #(18,FLUX) rd_add_18_40_opA(clk);
        read_interface #(18,FLUX) rd_add_18_40_opB(clk);
        write_interface #(18,FLUX) wr_add_18_40_sum(clk);

        //add_18_41
        read_interface #(18,FLUX) rd_add_18_41_opA(clk);
        read_interface #(18,FLUX) rd_add_18_41_opB(clk);
        write_interface #(18,FLUX) wr_add_18_41_sum(clk);

//7� riga               

        //add_18_42
        read_interface #(18,FLUX) rd_add_18_42_opA(clk);
        read_interface #(18,FLUX) rd_add_18_42_opB(clk);
        write_interface #(18,FLUX) wr_add_18_42_sum(clk);
        
        //add_18_43
        read_interface #(18,FLUX) rd_add_18_43_opA(clk);
        read_interface #(18,FLUX) rd_add_18_43_opB(clk);
        write_interface #(18,FLUX) wr_add_18_43_sum(clk);
        
        //add_18_44
        read_interface #(18,FLUX) rd_add_18_44_opA(clk);
        read_interface #(18,FLUX) rd_add_18_44_opB(clk);
        write_interface #(18,FLUX) wr_add_18_44_sum(clk);
        
        //add_18_45
        read_interface #(18,FLUX) rd_add_18_45_opA(clk);
        read_interface #(18,FLUX) rd_add_18_45_opB(clk);
        write_interface #(18,FLUX) wr_add_18_45_sum(clk);
        
        //add_18_46
        read_interface #(18,FLUX) rd_add_18_46_opA(clk);
        read_interface #(18,FLUX) rd_add_18_46_opB(clk);
        write_interface #(18,FLUX) wr_add_18_46_sum(clk);
        
        //add_18_47
        read_interface #(18,FLUX) rd_add_18_47_opA(clk);
        read_interface #(18,FLUX) rd_add_18_47_opB(clk);
        write_interface #(18,FLUX) wr_add_18_47_sum(clk);

        //add_18_48
        read_interface #(18,FLUX) rd_add_18_48_opA(clk);
        read_interface #(18,FLUX) rd_add_18_48_opB(clk);
        write_interface #(18,FLUX) wr_add_18_48_sum(clk);      
        
//8� riga               

        //add_18_49
        read_interface #(18,FLUX) rd_add_18_49_opA(clk);
        read_interface #(18,FLUX) rd_add_18_49_opB(clk);
        write_interface #(18,FLUX) wr_add_18_49_sum(clk);
        
        //add_18_50
        read_interface #(18,FLUX) rd_add_18_50_opA(clk);
        read_interface #(18,FLUX) rd_add_18_50_opB(clk);
        write_interface #(18,FLUX) wr_add_18_50_sum(clk);
        
        //add_18_51
        read_interface #(18,FLUX) rd_add_18_51_opA(clk);
        read_interface #(18,FLUX) rd_add_18_51_opB(clk);
        write_interface #(18,FLUX) wr_add_18_51_sum(clk);
        
        //add_18_52
        read_interface #(18,FLUX) rd_add_18_52_opA(clk);
        read_interface #(18,FLUX) rd_add_18_52_opB(clk);
        write_interface #(18,FLUX) wr_add_18_52_sum(clk);
        
        //add_18_53
        read_interface #(18,FLUX) rd_add_18_53_opA(clk);
        read_interface #(18,FLUX) rd_add_18_53_opB(clk);
        write_interface #(18,FLUX) wr_add_18_53_sum(clk);
        
        //add_18_54
        read_interface #(18,FLUX) rd_add_18_54_opA(clk);
        read_interface #(18,FLUX) rd_add_18_54_opB(clk);
        write_interface #(18,FLUX) wr_add_18_54_sum(clk);

        //add_18_55
        read_interface #(18,FLUX) rd_add_18_55_opA(clk);
        read_interface #(18,FLUX) rd_add_18_55_opB(clk);
        write_interface #(18,FLUX) wr_add_18_55_sum(clk);                         

    //COEFF LUMA H

        //coeff_luma_h
        read_interface #(3,FLUX) rd_coeff_luma_h_alpha(clk);
        write_interface #(9,FLUX) wr_coeff_luma_h_c0(clk);
        write_interface #(9,FLUX) wr_coeff_luma_h_c1(clk);
        write_interface #(9,FLUX) wr_coeff_luma_h_c2(clk);
        write_interface #(9,FLUX) wr_coeff_luma_h_c3(clk);
        write_interface #(9,FLUX) wr_coeff_luma_h_c4(clk);
        write_interface #(9,FLUX) wr_coeff_luma_h_c5(clk);
        write_interface #(9,FLUX) wr_coeff_luma_h_c6(clk);
        write_interface #(9,FLUX) wr_coeff_luma_h_c7(clk);

    //DERIVE REAL SIZE (x1)
        
        //derive_real_size
        read_interface #(7,FLUX) rd_derive_real_size_ext_size(clk);
        write_interface #(7,FLUX) wr_derive_real_size_real_size(clk);

    //REMOVE H (x1)
    
        //remove_h
        read_interface #(7,FLUX) rd_remove_h_0_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_h_1_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_h_2_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_h_3_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_h_4_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_h_5_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_h_6_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_h_7_ext_size(clk);
        read_interface #(18,FLUX) rd_remove_h_0_in_pel(clk);
        read_interface #(18,FLUX) rd_remove_h_1_in_pel(clk);
        read_interface #(18,FLUX) rd_remove_h_2_in_pel(clk);
        read_interface #(18,FLUX) rd_remove_h_3_in_pel(clk);
        read_interface #(18,FLUX) rd_remove_h_4_in_pel(clk);
        read_interface #(18,FLUX) rd_remove_h_5_in_pel(clk);
        read_interface #(18,FLUX) rd_remove_h_6_in_pel(clk);
        read_interface #(18,FLUX) rd_remove_h_7_in_pel(clk);                            
        write_interface #(18,FLUX) wr_remove_h_0_out_pel(clk);
        write_interface #(18,FLUX) wr_remove_h_1_out_pel(clk);
        write_interface #(18,FLUX) wr_remove_h_2_out_pel(clk);
        write_interface #(18,FLUX) wr_remove_h_3_out_pel(clk);
        write_interface #(18,FLUX) wr_remove_h_4_out_pel(clk);
        write_interface #(18,FLUX) wr_remove_h_5_out_pel(clk);
        write_interface #(18,FLUX) wr_remove_h_6_out_pel(clk);
        write_interface #(18,FLUX) wr_remove_h_7_out_pel(clk);
                        
//SECONDA PARTE

    //REMOVE V (x1)
    
        //remove_v
        read_interface #(7,FLUX) rd_remove_v_0_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_v_1_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_v_2_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_v_3_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_v_4_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_v_5_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_v_6_ext_size(clk);
		read_interface #(7,FLUX) rd_remove_v_7_ext_size(clk);
        read_interface #(7,FLUX) rd_remove_v_0_real_size(clk);
		read_interface #(7,FLUX) rd_remove_v_1_real_size(clk);
		read_interface #(7,FLUX) rd_remove_v_2_real_size(clk);
		read_interface #(7,FLUX) rd_remove_v_3_real_size(clk);
		read_interface #(7,FLUX) rd_remove_v_4_real_size(clk);
		read_interface #(7,FLUX) rd_remove_v_5_real_size(clk);
		read_interface #(7,FLUX) rd_remove_v_6_real_size(clk);
		read_interface #(7,FLUX) rd_remove_v_7_real_size(clk);
        read_interface #(8,FLUX) rd_remove_v_0_in_pel(clk);
        read_interface #(8,FLUX) rd_remove_v_1_in_pel(clk);
        read_interface #(8,FLUX) rd_remove_v_2_in_pel(clk);
        read_interface #(8,FLUX) rd_remove_v_3_in_pel(clk);
        read_interface #(8,FLUX) rd_remove_v_4_in_pel(clk);
        read_interface #(8,FLUX) rd_remove_v_5_in_pel(clk);
        read_interface #(8,FLUX) rd_remove_v_6_in_pel(clk);
        read_interface #(8,FLUX) rd_remove_v_7_in_pel(clk);    
        write_interface #(8,FLUX) wr_remove_v_0_out_pel(clk);
        write_interface #(8,FLUX) wr_remove_v_1_out_pel(clk);
        write_interface #(8,FLUX) wr_remove_v_2_out_pel(clk);
        write_interface #(8,FLUX) wr_remove_v_3_out_pel(clk);
        write_interface #(8,FLUX) wr_remove_v_4_out_pel(clk);
        write_interface #(8,FLUX) wr_remove_v_5_out_pel(clk);
        write_interface #(8,FLUX) wr_remove_v_6_out_pel(clk);
        write_interface #(8,FLUX) wr_remove_v_7_out_pel(clk);

    //CLIP (x8)
    
        //clip_0
        read_interface #(16,FLUX) rd_clip_0_in_pel(clk);
        write_interface #(8,FLUX) wr_clip_0_out_pel(clk);

        //clip_1
        read_interface #(16,FLUX) rd_clip_1_in_pel(clk);
        write_interface #(8,FLUX) wr_clip_1_out_pel(clk);
        
        //clip_2
        read_interface #(16,FLUX) rd_clip_2_in_pel(clk);
        write_interface #(8,FLUX) wr_clip_2_out_pel(clk);
        
        //clip_3
        read_interface #(16,FLUX) rd_clip_3_in_pel(clk);
        write_interface #(8,FLUX) wr_clip_3_out_pel(clk);

        //clip_4
        read_interface #(16,FLUX) rd_clip_4_in_pel(clk);
        write_interface #(8,FLUX) wr_clip_4_out_pel(clk);
        
        //clip_5
        read_interface #(16,FLUX) rd_clip_5_in_pel(clk);
        write_interface #(8,FLUX) wr_clip_5_out_pel(clk);

        //clip_6
        read_interface #(16,FLUX) rd_clip_6_in_pel(clk);
        write_interface #(8,FLUX) wr_clip_6_out_pel(clk);
        
        //clip_7
        read_interface #(16,FLUX) rd_clip_7_in_pel(clk);
        write_interface #(8,FLUX) wr_clip_7_out_pel(clk);                            
            
    //SHIFT (x8)
    
        //shift_0
        read_interface #(27,FLUX) rd_shift_0_in_pel(clk);
        write_interface #(16,FLUX) wr_shift_0_out_pel(clk);

        //shift_1
        read_interface #(27,FLUX) rd_shift_1_in_pel(clk);
        write_interface #(16,FLUX) wr_shift_1_out_pel(clk);        

        //shift_2
        read_interface #(27,FLUX) rd_shift_2_in_pel(clk);
        write_interface #(16,FLUX) wr_shift_2_out_pel(clk);

        //shift_3
        read_interface #(27,FLUX) rd_shift_3_in_pel(clk);
        write_interface #(16,FLUX) wr_shift_3_out_pel(clk);

        //shift_4
        read_interface #(27,FLUX) rd_shift_4_in_pel(clk);
        write_interface #(16,FLUX) wr_shift_4_out_pel(clk);

        //shift_5
        read_interface #(27,FLUX) rd_shift_5_in_pel(clk);
        write_interface #(16,FLUX) wr_shift_5_out_pel(clk);        

        //shift_6
        read_interface #(27,FLUX) rd_shift_6_in_pel(clk);
        write_interface #(16,FLUX) wr_shift_6_out_pel(clk);

        //shift_7
        read_interface #(27,FLUX) rd_shift_7_in_pel(clk);
        write_interface #(16,FLUX) wr_shift_7_out_pel(clk);        

    //COEFF LUMA V (x1)

        //coeff_luma_v
        read_interface #(3,FLUX) rd_coeff_luma_v_alpha(clk);
        write_interface #(9,FLUX) wr_coeff_luma_v_c0(clk);
        write_interface #(9,FLUX) wr_coeff_luma_v_c1(clk);
        write_interface #(9,FLUX) wr_coeff_luma_v_c2(clk);
        write_interface #(9,FLUX) wr_coeff_luma_v_c3(clk);
        write_interface #(9,FLUX) wr_coeff_luma_v_c4(clk);
        write_interface #(9,FLUX) wr_coeff_luma_v_c5(clk);
        write_interface #(9,FLUX) wr_coeff_luma_v_c6(clk);
        write_interface #(9,FLUX) wr_coeff_luma_v_c7(clk);

    //LINE BUFFER (x7)
    
        //line_buffer_0
        read_interface #(7,FLUX) rd_line_buffer_0_real_size(clk);
        read_interface #(7,FLUX) rd_line_buffer_0_ext_size(clk);
        read_interface #(18,FLUX) rd_line_buffer_0_0_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_0_1_in_pel(clk);        
        read_interface #(18,FLUX) rd_line_buffer_0_2_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_0_3_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_0_4_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_0_5_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_0_6_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_0_7_in_pel(clk);                                                    
        write_interface #(18,FLUX) wr_line_buffer_0_0_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_0_1_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_0_2_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_0_3_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_0_4_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_0_5_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_0_6_out_pel(clk);                        
        write_interface #(18,FLUX) wr_line_buffer_0_7_out_pel(clk);                                
    
        //line_buffer_1
        read_interface #(7,FLUX) rd_line_buffer_1_real_size(clk);
        read_interface #(7,FLUX) rd_line_buffer_1_ext_size(clk);
        read_interface #(18,FLUX) rd_line_buffer_1_0_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_1_1_in_pel(clk);        
        read_interface #(18,FLUX) rd_line_buffer_1_2_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_1_3_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_1_4_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_1_5_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_1_6_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_1_7_in_pel(clk);                                                    
        write_interface #(18,FLUX) wr_line_buffer_1_0_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_1_1_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_1_2_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_1_3_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_1_4_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_1_5_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_1_6_out_pel(clk);                        
        write_interface #(18,FLUX) wr_line_buffer_1_7_out_pel(clk);
    
        //line_buffer_2
        read_interface #(7,FLUX) rd_line_buffer_2_real_size(clk);
        read_interface #(7,FLUX) rd_line_buffer_2_ext_size(clk);
        read_interface #(18,FLUX) rd_line_buffer_2_0_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_2_1_in_pel(clk);        
        read_interface #(18,FLUX) rd_line_buffer_2_2_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_2_3_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_2_4_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_2_5_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_2_6_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_2_7_in_pel(clk);                                                    
        write_interface #(18,FLUX) wr_line_buffer_2_0_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_2_1_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_2_2_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_2_3_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_2_4_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_2_5_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_2_6_out_pel(clk);                        
        write_interface #(18,FLUX) wr_line_buffer_2_7_out_pel(clk);
        
        //line_buffer_3
        read_interface #(7,FLUX) rd_line_buffer_3_real_size(clk);
        read_interface #(7,FLUX) rd_line_buffer_3_ext_size(clk);
        read_interface #(18,FLUX) rd_line_buffer_3_0_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_3_1_in_pel(clk);        
        read_interface #(18,FLUX) rd_line_buffer_3_2_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_3_3_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_3_4_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_3_5_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_3_6_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_3_7_in_pel(clk);                                                    
        write_interface #(18,FLUX) wr_line_buffer_3_0_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_3_1_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_3_2_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_3_3_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_3_4_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_3_5_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_3_6_out_pel(clk);                        
        write_interface #(18,FLUX) wr_line_buffer_3_7_out_pel(clk);
        
        //line_buffer_4
        read_interface #(7,FLUX) rd_line_buffer_4_real_size(clk);
        read_interface #(7,FLUX) rd_line_buffer_4_ext_size(clk);
        read_interface #(18,FLUX) rd_line_buffer_4_0_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_4_1_in_pel(clk);        
        read_interface #(18,FLUX) rd_line_buffer_4_2_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_4_3_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_4_4_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_4_5_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_4_6_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_4_7_in_pel(clk);                                                    
        write_interface #(18,FLUX) wr_line_buffer_4_0_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_4_1_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_4_2_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_4_3_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_4_4_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_4_5_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_4_6_out_pel(clk);                        
        write_interface #(18,FLUX) wr_line_buffer_4_7_out_pel(clk);
        
        //line_buffer_5
        read_interface #(7,FLUX) rd_line_buffer_5_real_size(clk);
        read_interface #(7,FLUX) rd_line_buffer_5_ext_size(clk);
        read_interface #(18,FLUX) rd_line_buffer_5_0_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_5_1_in_pel(clk);        
        read_interface #(18,FLUX) rd_line_buffer_5_2_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_5_3_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_5_4_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_5_5_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_5_6_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_5_7_in_pel(clk);                                                    
        write_interface #(18,FLUX) wr_line_buffer_5_0_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_5_1_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_5_2_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_5_3_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_5_4_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_5_5_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_5_6_out_pel(clk);                        
        write_interface #(18,FLUX) wr_line_buffer_5_7_out_pel(clk);
    
        //line_buffer_6
        read_interface #(7,FLUX) rd_line_buffer_6_real_size(clk);
        read_interface #(7,FLUX) rd_line_buffer_6_ext_size(clk);
        read_interface #(18,FLUX) rd_line_buffer_6_0_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_6_1_in_pel(clk);        
        read_interface #(18,FLUX) rd_line_buffer_6_2_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_6_3_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_6_4_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_6_5_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_6_6_in_pel(clk);
        read_interface #(18,FLUX) rd_line_buffer_6_7_in_pel(clk);                                                    
        write_interface #(18,FLUX) wr_line_buffer_6_0_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_6_1_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_6_2_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_6_3_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_6_4_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_6_5_out_pel(clk);
        write_interface #(18,FLUX) wr_line_buffer_6_6_out_pel(clk);                        
        write_interface #(18,FLUX) wr_line_buffer_6_7_out_pel(clk);

        
    //MUL_18 (x64)        
        
//1�colonna
    
        //mul_18_0
        read_interface #(7,FLUX) rd_mul_18_0_real_size(clk);
        read_interface #(7,FLUX) rd_mul_18_0_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_0_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_0_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_0_prod(clk);
        
        //mul_18_1
        read_interface #(7,FLUX) rd_mul_18_1_real_size(clk);
        read_interface #(7,FLUX) rd_mul_18_1_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_1_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_1_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_1_prod(clk);
        
        //mul_18_2
        read_interface #(7,FLUX) rd_mul_18_2_real_size(clk);
        read_interface #(7,FLUX) rd_mul_18_2_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_2_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_2_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_2_prod(clk);
                
        //mul_18_3
        read_interface #(7,FLUX) rd_mul_18_3_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_3_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_3_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_3_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_3_prod(clk);
        
        //mul_18_4
        read_interface #(7,FLUX) rd_mul_18_4_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_4_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_4_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_4_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_4_prod(clk);
        
        //mul_18_5
        read_interface #(7,FLUX) rd_mul_18_5_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_5_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_5_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_5_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_5_prod(clk);
        
        //mul_18_6
        read_interface #(7,FLUX) rd_mul_18_6_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_6_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_6_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_6_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_6_prod(clk);
                
        //mul_18_7
        read_interface #(7,FLUX) rd_mul_18_7_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_7_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_7_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_7_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_7_prod(clk);

//2�colonna
    
        //mul_18_8
        read_interface #(7,FLUX) rd_mul_18_8_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_8_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_8_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_8_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_8_prod(clk);
        
        //mul_18_9
        read_interface #(7,FLUX) rd_mul_18_9_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_9_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_9_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_9_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_9_prod(clk);
        
        //mul_18_10
        read_interface #(7,FLUX) rd_mul_18_10_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_10_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_10_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_10_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_10_prod(clk);
                
        //mul_18_11
        read_interface #(7,FLUX) rd_mul_18_11_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_11_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_11_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_11_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_11_prod(clk);
        
        //mul_18_12
        read_interface #(7,FLUX) rd_mul_18_12_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_12_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_12_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_12_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_12_prod(clk);
        
        //mul_18_13
        read_interface #(7,FLUX) rd_mul_18_13_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_13_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_13_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_13_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_13_prod(clk);
        
        //mul_18_14
        read_interface #(7,FLUX) rd_mul_18_14_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_14_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_14_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_14_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_14_prod(clk);
                
        //mul_18_15
        read_interface #(7,FLUX) rd_mul_18_15_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_15_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_15_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_15_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_15_prod(clk);

//3�colonna
    
        //mul_18_16
        read_interface #(7,FLUX) rd_mul_18_16_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_16_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_16_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_16_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_16_prod(clk);
        
        //mul_18_17
        read_interface #(7,FLUX) rd_mul_18_17_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_17_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_17_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_17_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_17_prod(clk);
        
        //mul_18_18
        read_interface #(7,FLUX) rd_mul_18_18_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_18_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_18_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_18_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_18_prod(clk);
                
        //mul_18_19
        read_interface #(7,FLUX) rd_mul_18_19_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_19_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_19_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_19_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_19_prod(clk);
        
        //mul_18_20
        read_interface #(7,FLUX) rd_mul_18_20_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_20_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_20_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_20_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_20_prod(clk);
        
        //mul_18_21
        read_interface #(7,FLUX) rd_mul_18_21_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_21_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_21_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_21_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_21_prod(clk);
        
        //mul_18_22
        read_interface #(7,FLUX) rd_mul_18_22_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_22_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_22_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_22_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_22_prod(clk);
                
        //mul_18_23
        read_interface #(7,FLUX) rd_mul_18_23_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_23_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_23_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_23_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_23_prod(clk);

//4�colonna
    
        //mul_18_24
        read_interface #(7,FLUX) rd_mul_18_24_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_24_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_24_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_24_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_24_prod(clk);
        
        //mul_18_25
        read_interface #(7,FLUX) rd_mul_18_25_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_25_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_25_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_25_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_25_prod(clk);
        
        //mul_18_26
        read_interface #(7,FLUX) rd_mul_18_26_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_26_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_26_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_26_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_26_prod(clk);
                
        //mul_18_27
        read_interface #(7,FLUX) rd_mul_18_27_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_27_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_27_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_27_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_27_prod(clk);
        
        //mul_18_28
        read_interface #(7,FLUX) rd_mul_18_28_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_28_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_28_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_28_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_28_prod(clk);
        
        //mul_18_29
        read_interface #(7,FLUX) rd_mul_18_29_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_29_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_29_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_29_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_29_prod(clk);
        
        //mul_18_30
        read_interface #(7,FLUX) rd_mul_18_30_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_30_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_30_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_30_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_30_prod(clk);
                
        //mul_18_31
        read_interface #(7,FLUX) rd_mul_18_31_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_31_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_31_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_31_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_31_prod(clk);

//5�colonna
    
        //mul_18_32
        read_interface #(7,FLUX) rd_mul_18_32_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_32_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_32_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_32_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_32_prod(clk);
        
        //mul_18_33
        read_interface #(7,FLUX) rd_mul_18_33_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_33_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_33_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_33_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_33_prod(clk);
        
        //mul_18_34
        read_interface #(7,FLUX) rd_mul_18_34_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_34_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_34_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_34_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_34_prod(clk);
                
        //mul_18_35
        read_interface #(7,FLUX) rd_mul_18_35_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_35_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_35_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_35_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_35_prod(clk);
        
        //mul_18_36
        read_interface #(7,FLUX) rd_mul_18_36_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_36_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_36_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_36_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_36_prod(clk);
        
        //mul_18_37
        read_interface #(7,FLUX) rd_mul_18_37_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_37_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_37_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_37_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_37_prod(clk);
        
        //mul_18_38
        read_interface #(7,FLUX) rd_mul_18_38_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_38_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_38_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_38_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_38_prod(clk);
                
        //mul_18_39
        read_interface #(7,FLUX) rd_mul_18_39_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_39_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_39_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_39_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_39_prod(clk);

//6�colonna
    
        //mul_18_40
        read_interface #(7,FLUX) rd_mul_18_40_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_40_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_40_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_40_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_40_prod(clk);
        
        //mul_18_41
        read_interface #(7,FLUX) rd_mul_18_41_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_41_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_41_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_41_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_41_prod(clk);
        
        //mul_18_42
        read_interface #(7,FLUX) rd_mul_18_42_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_42_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_42_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_42_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_42_prod(clk);
                
        //mul_18_43
        read_interface #(7,FLUX) rd_mul_18_43_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_43_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_43_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_43_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_43_prod(clk);
        
        //mul_18_44
        read_interface #(7,FLUX) rd_mul_18_44_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_44_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_44_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_44_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_44_prod(clk);
        
        //mul_18_45
        read_interface #(7,FLUX) rd_mul_18_45_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_45_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_45_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_45_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_45_prod(clk);
        
        //mul_18_46
        read_interface #(7,FLUX) rd_mul_18_46_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_46_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_46_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_46_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_46_prod(clk);
                
        //mul_18_47
        read_interface #(7,FLUX) rd_mul_18_47_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_47_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_47_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_47_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_47_prod(clk);
        

//7�colonna
    
        //mul_18_48
        read_interface #(7,FLUX) rd_mul_18_48_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_48_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_48_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_48_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_48_prod(clk);
        
        //mul_18_49
        read_interface #(7,FLUX) rd_mul_18_49_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_49_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_49_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_49_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_49_prod(clk);
        
        //mul_18_50
        read_interface #(7,FLUX) rd_mul_18_50_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_50_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_50_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_50_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_50_prod(clk);
                
        //mul_18_51
        read_interface #(7,FLUX) rd_mul_18_51_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_51_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_51_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_51_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_51_prod(clk);
        
        //mul_18_52
        read_interface #(7,FLUX) rd_mul_18_52_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_52_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_52_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_52_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_52_prod(clk);
        
        //mul_18_53
        read_interface #(7,FLUX) rd_mul_18_53_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_53_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_53_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_53_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_53_prod(clk);
        
        //mul_18_54
        read_interface #(7,FLUX) rd_mul_18_54_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_54_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_54_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_54_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_54_prod(clk);
                
        //mul_18_55
        read_interface #(7,FLUX) rd_mul_18_55_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_55_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_55_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_55_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_55_prod(clk);        


//8�colonna
    
        //mul_18_56
        read_interface #(7,FLUX) rd_mul_18_56_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_56_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_56_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_56_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_56_prod(clk);
        
        //mul_18_57
        read_interface #(7,FLUX) rd_mul_18_57_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_57_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_57_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_57_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_57_prod(clk);
        
        //mul_18_58
        read_interface #(7,FLUX) rd_mul_18_58_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_58_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_58_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_58_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_58_prod(clk);
                
        //mul_18_59
        read_interface #(7,FLUX) rd_mul_18_59_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_59_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_59_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_59_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_59_prod(clk);
        
        //mul_18_60
        read_interface #(7,FLUX) rd_mul_18_60_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_60_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_60_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_60_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_60_prod(clk);
        
        //mul_18_61
        read_interface #(7,FLUX) rd_mul_18_61_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_61_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_61_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_61_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_61_prod(clk);
        
        //mul_18_62
        read_interface #(7,FLUX) rd_mul_18_62_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_62_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_62_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_62_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_62_prod(clk);
                
        //mul_18_63
        read_interface #(7,FLUX) rd_mul_18_63_real_size(clk);        
        read_interface #(7,FLUX) rd_mul_18_63_ext_size(clk);
        read_interface #(18,FLUX) rd_mul_18_63_opA(clk);
        read_interface #(9,FLUX) rd_mul_18_63_opB(clk);
        write_interface #(27,FLUX) wr_mul_18_63_prod(clk);
    
    //ADD_27 (x56) 

//1� riga
    
        //add_27_0
        read_interface #(27,FLUX) rd_add_27_0_opA(clk);
        read_interface #(27,FLUX) rd_add_27_0_opB(clk);
        write_interface #(27,FLUX) wr_add_27_0_sum(clk);
        
        //add_27_1
        read_interface #(27,FLUX) rd_add_27_1_opA(clk);
        read_interface #(27,FLUX) rd_add_27_1_opB(clk);
        write_interface #(27,FLUX) wr_add_27_1_sum(clk);
        
        //add_27_2
        read_interface #(27,FLUX) rd_add_27_2_opA(clk);
        read_interface #(27,FLUX) rd_add_27_2_opB(clk);
        write_interface #(27,FLUX) wr_add_27_2_sum(clk);
        
        //add_27_3
        read_interface #(27,FLUX) rd_add_27_3_opA(clk);
        read_interface #(27,FLUX) rd_add_27_3_opB(clk);
        write_interface #(27,FLUX) wr_add_27_3_sum(clk);
        
        //add_27_4
        read_interface #(27,FLUX) rd_add_27_4_opA(clk);
        read_interface #(27,FLUX) rd_add_27_4_opB(clk);
        write_interface #(27,FLUX) wr_add_27_4_sum(clk);
        
        //add_27_5
        read_interface #(27,FLUX) rd_add_27_5_opA(clk);
        read_interface #(27,FLUX) rd_add_27_5_opB(clk);
        write_interface #(27,FLUX) wr_add_27_5_sum(clk);

        //add_27_6
        read_interface #(27,FLUX) rd_add_27_6_opA(clk);
        read_interface #(27,FLUX) rd_add_27_6_opB(clk);
        write_interface #(27,FLUX) wr_add_27_6_sum(clk);        

//2� riga
    
        //add_27_7
        read_interface #(27,FLUX) rd_add_27_7_opA(clk);
        read_interface #(27,FLUX) rd_add_27_7_opB(clk);
        write_interface #(27,FLUX) wr_add_27_7_sum(clk);
        
        //add_27_8
        read_interface #(27,FLUX) rd_add_27_8_opA(clk);
        read_interface #(27,FLUX) rd_add_27_8_opB(clk);
        write_interface #(27,FLUX) wr_add_27_8_sum(clk);
        
        //add_27_9
        read_interface #(27,FLUX) rd_add_27_9_opA(clk);
        read_interface #(27,FLUX) rd_add_27_9_opB(clk);
        write_interface #(27,FLUX) wr_add_27_9_sum(clk);
        
        //add_27_10
        read_interface #(27,FLUX) rd_add_27_10_opA(clk);
        read_interface #(27,FLUX) rd_add_27_10_opB(clk);
        write_interface #(27,FLUX) wr_add_27_10_sum(clk);
        
        //add_27_11
        read_interface #(27,FLUX) rd_add_27_11_opA(clk);
        read_interface #(27,FLUX) rd_add_27_11_opB(clk);
        write_interface #(27,FLUX) wr_add_27_11_sum(clk);
        
        //add_27_12
        read_interface #(27,FLUX) rd_add_27_12_opA(clk);
        read_interface #(27,FLUX) rd_add_27_12_opB(clk);
        write_interface #(27,FLUX) wr_add_27_12_sum(clk);

        //add_27_13
        read_interface #(27,FLUX) rd_add_27_13_opA(clk);
        read_interface #(27,FLUX) rd_add_27_13_opB(clk);
        write_interface #(27,FLUX) wr_add_27_13_sum(clk);
        
//3� riga
    
        //add_27_14
        read_interface #(27,FLUX) rd_add_27_14_opA(clk);
        read_interface #(27,FLUX) rd_add_27_14_opB(clk);
        write_interface #(27,FLUX) wr_add_27_14_sum(clk);
        
        //add_27_15
        read_interface #(27,FLUX) rd_add_27_15_opA(clk);
        read_interface #(27,FLUX) rd_add_27_15_opB(clk);
        write_interface #(27,FLUX) wr_add_27_15_sum(clk);
        
        //add_27_16
        read_interface #(27,FLUX) rd_add_27_16_opA(clk);
        read_interface #(27,FLUX) rd_add_27_16_opB(clk);
        write_interface #(27,FLUX) wr_add_27_16_sum(clk);
        
        //add_27_17
        read_interface #(27,FLUX) rd_add_27_17_opA(clk);
        read_interface #(27,FLUX) rd_add_27_17_opB(clk);
        write_interface #(27,FLUX) wr_add_27_17_sum(clk);
        
        //add_27_18
        read_interface #(27,FLUX) rd_add_27_18_opA(clk);
        read_interface #(27,FLUX) rd_add_27_18_opB(clk);
        write_interface #(27,FLUX) wr_add_27_18_sum(clk);
        
        //add_27_19
        read_interface #(27,FLUX) rd_add_27_19_opA(clk);
        read_interface #(27,FLUX) rd_add_27_19_opB(clk);
        write_interface #(27,FLUX) wr_add_27_19_sum(clk);

        //add_27_20
        read_interface #(27,FLUX) rd_add_27_20_opA(clk);
        read_interface #(27,FLUX) rd_add_27_20_opB(clk);
        write_interface #(27,FLUX) wr_add_27_20_sum(clk);                 
        
//4� riga
    
        //add_27_21
        read_interface #(27,FLUX) rd_add_27_21_opA(clk);
        read_interface #(27,FLUX) rd_add_27_21_opB(clk);
        write_interface #(27,FLUX) wr_add_27_21_sum(clk);
        
        //add_27_22
        read_interface #(27,FLUX) rd_add_27_22_opA(clk);
        read_interface #(27,FLUX) rd_add_27_22_opB(clk);
        write_interface #(27,FLUX) wr_add_27_22_sum(clk);
        
        //add_27_23
        read_interface #(27,FLUX) rd_add_27_23_opA(clk);
        read_interface #(27,FLUX) rd_add_27_23_opB(clk);
        write_interface #(27,FLUX) wr_add_27_23_sum(clk);
        
        //add_27_24
        read_interface #(27,FLUX) rd_add_27_24_opA(clk);
        read_interface #(27,FLUX) rd_add_27_24_opB(clk);
        write_interface #(27,FLUX) wr_add_27_24_sum(clk);
        
        //add_27_25
        read_interface #(27,FLUX) rd_add_27_25_opA(clk);
        read_interface #(27,FLUX) rd_add_27_25_opB(clk);
        write_interface #(27,FLUX) wr_add_27_25_sum(clk);
        
        //add_27_26
        read_interface #(27,FLUX) rd_add_27_26_opA(clk);
        read_interface #(27,FLUX) rd_add_27_26_opB(clk);
        write_interface #(27,FLUX) wr_add_27_26_sum(clk);

        //add_27_27
        read_interface #(27,FLUX) rd_add_27_27_opA(clk);
        read_interface #(27,FLUX) rd_add_27_27_opB(clk);
        write_interface #(27,FLUX) wr_add_27_27_sum(clk); 
        
//5� riga               

        //add_27_28
        read_interface #(27,FLUX) rd_add_27_28_opA(clk);
        read_interface #(27,FLUX) rd_add_27_28_opB(clk);
        write_interface #(27,FLUX) wr_add_27_28_sum(clk);
        
        //add_27_29
        read_interface #(27,FLUX) rd_add_27_29_opA(clk);
        read_interface #(27,FLUX) rd_add_27_29_opB(clk);
        write_interface #(27,FLUX) wr_add_27_29_sum(clk);
        
        //add_27_30
        read_interface #(27,FLUX) rd_add_27_30_opA(clk);
        read_interface #(27,FLUX) rd_add_27_30_opB(clk);
        write_interface #(27,FLUX) wr_add_27_30_sum(clk);
        
        //add_27_31
        read_interface #(27,FLUX) rd_add_27_31_opA(clk);
        read_interface #(27,FLUX) rd_add_27_31_opB(clk);
        write_interface #(27,FLUX) wr_add_27_31_sum(clk);
        
        //add_27_32
        read_interface #(27,FLUX) rd_add_27_32_opA(clk);
        read_interface #(27,FLUX) rd_add_27_32_opB(clk);
        write_interface #(27,FLUX) wr_add_27_32_sum(clk);
        
        //add_27_33
        read_interface #(27,FLUX) rd_add_27_33_opA(clk);
        read_interface #(27,FLUX) rd_add_27_33_opB(clk);
        write_interface #(27,FLUX) wr_add_27_33_sum(clk);

        //add_27_34
        read_interface #(27,FLUX) rd_add_27_34_opA(clk);
        read_interface #(27,FLUX) rd_add_27_34_opB(clk);
        write_interface #(27,FLUX) wr_add_27_34_sum(clk);

//6� riga               

        //add_27_35
        read_interface #(27,FLUX) rd_add_27_35_opA(clk);
        read_interface #(27,FLUX) rd_add_27_35_opB(clk);
        write_interface #(27,FLUX) wr_add_27_35_sum(clk);
        
        //add_27_36
        read_interface #(27,FLUX) rd_add_27_36_opA(clk);
        read_interface #(27,FLUX) rd_add_27_36_opB(clk);
        write_interface #(27,FLUX) wr_add_27_36_sum(clk);
        
        //add_27_37
        read_interface #(27,FLUX) rd_add_27_37_opA(clk);
        read_interface #(27,FLUX) rd_add_27_37_opB(clk);
        write_interface #(27,FLUX) wr_add_27_37_sum(clk);
        
        //add_27_38
        read_interface #(27,FLUX) rd_add_27_38_opA(clk);
        read_interface #(27,FLUX) rd_add_27_38_opB(clk);
        write_interface #(27,FLUX) wr_add_27_38_sum(clk);
        
        //add_27_39
        read_interface #(27,FLUX) rd_add_27_39_opA(clk);
        read_interface #(27,FLUX) rd_add_27_39_opB(clk);
        write_interface #(27,FLUX) wr_add_27_39_sum(clk);
        
        //add_27_40
        read_interface #(27,FLUX) rd_add_27_40_opA(clk);
        read_interface #(27,FLUX) rd_add_27_40_opB(clk);
        write_interface #(27,FLUX) wr_add_27_40_sum(clk);

        //add_27_41
        read_interface #(27,FLUX) rd_add_27_41_opA(clk);
        read_interface #(27,FLUX) rd_add_27_41_opB(clk);
        write_interface #(27,FLUX) wr_add_27_41_sum(clk);

//7� riga               

        //add_27_42
        read_interface #(27,FLUX) rd_add_27_42_opA(clk);
        read_interface #(27,FLUX) rd_add_27_42_opB(clk);
        write_interface #(27,FLUX) wr_add_27_42_sum(clk);
        
        //add_27_43
        read_interface #(27,FLUX) rd_add_27_43_opA(clk);
        read_interface #(27,FLUX) rd_add_27_43_opB(clk);
        write_interface #(27,FLUX) wr_add_27_43_sum(clk);
        
        //add_27_44
        read_interface #(27,FLUX) rd_add_27_44_opA(clk);
        read_interface #(27,FLUX) rd_add_27_44_opB(clk);
        write_interface #(27,FLUX) wr_add_27_44_sum(clk);
        
        //add_27_45
        read_interface #(27,FLUX) rd_add_27_45_opA(clk);
        read_interface #(27,FLUX) rd_add_27_45_opB(clk);
        write_interface #(27,FLUX) wr_add_27_45_sum(clk);
        
        //add_27_46
        read_interface #(27,FLUX) rd_add_27_46_opA(clk);
        read_interface #(27,FLUX) rd_add_27_46_opB(clk);
        write_interface #(27,FLUX) wr_add_27_46_sum(clk);
        
        //add_27_47
        read_interface #(27,FLUX) rd_add_27_47_opA(clk);
        read_interface #(27,FLUX) rd_add_27_47_opB(clk);
        write_interface #(27,FLUX) wr_add_27_47_sum(clk);

        //add_27_48
        read_interface #(27,FLUX) rd_add_27_48_opA(clk);
        read_interface #(27,FLUX) rd_add_27_48_opB(clk);
        write_interface #(27,FLUX) wr_add_27_48_sum(clk);      
        
//8� riga               

        //add_27_49
        read_interface #(27,FLUX) rd_add_27_49_opA(clk);
        read_interface #(27,FLUX) rd_add_27_49_opB(clk);
        write_interface #(27,FLUX) wr_add_27_49_sum(clk);
        
        //add_27_50
        read_interface #(27,FLUX) rd_add_27_50_opA(clk);
        read_interface #(27,FLUX) rd_add_27_50_opB(clk);
        write_interface #(27,FLUX) wr_add_27_50_sum(clk);
        
        //add_27_51
        read_interface #(27,FLUX) rd_add_27_51_opA(clk);
        read_interface #(27,FLUX) rd_add_27_51_opB(clk);
        write_interface #(27,FLUX) wr_add_27_51_sum(clk);
        
        //add_27_52
        read_interface #(27,FLUX) rd_add_27_52_opA(clk);
        read_interface #(27,FLUX) rd_add_27_52_opB(clk);
        write_interface #(27,FLUX) wr_add_27_52_sum(clk);
        
        //add_27_53
        read_interface #(27,FLUX) rd_add_27_53_opA(clk);
        read_interface #(27,FLUX) rd_add_27_53_opB(clk);
        write_interface #(27,FLUX) wr_add_27_53_sum(clk);
        
        //add_27_54
        read_interface #(27,FLUX) rd_add_27_54_opA(clk);
        read_interface #(27,FLUX) rd_add_27_54_opB(clk);
        write_interface #(27,FLUX) wr_add_27_54_sum(clk);

        //add_27_55
        read_interface #(27,FLUX) rd_add_27_55_opA(clk);
        read_interface #(27,FLUX) rd_add_27_55_opB(clk);
        write_interface #(27,FLUX) wr_add_27_55_sum(clk);                         



//FINE INTERFACCE MODULI




//FORKS



    //FORK MUL_9_0 / MUL_9_1 / MUL_9_2 / MUL_9_3 / MUL_9_4 / MUL_9_5 / MUL_9_6 / ... / MUL_9_63 / REMOVE_H ...
    //... / MUL_18_0 / MUL_18_1 / MUL_18_2 / MUL_18_3 / MUL_18_4 / MUL_18_5 / MUL_18_6 / ... / MUL_18_63 ...
    //... / REMOVE_v / LINE_BUFFER_0 / LINE_BUFFER_1 / LINE_BUFFER_2 / LINE_BUFFER_3 / LINE_BUFFER_4 ...
    //... / LINE_BUFFER_5 / LINE_BUFFER_6  / DERIVE_REAL_SIZE...
    //... ON EXTSIZE 
        
        // - INTERFACES
        
            //MUL9 (x64)
            
            //1� riga
            write_interface #(7,FLUX) wr_fifo_mul_9_0_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_1_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_2_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_3_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_4_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_5_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_6_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_7_ext_size (clk);
            //2� riga
            write_interface #(7,FLUX) wr_fifo_mul_9_8_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_9_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_10_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_11_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_12_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_13_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_14_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_15_ext_size (clk);            
            //3� riga
            write_interface #(7,FLUX) wr_fifo_mul_9_16_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_17_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_18_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_19_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_20_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_21_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_22_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_23_ext_size (clk);
            //4� riga
            write_interface #(7,FLUX) wr_fifo_mul_9_24_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_25_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_26_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_27_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_28_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_29_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_30_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_31_ext_size (clk);
            //5� riga
            write_interface #(7,FLUX) wr_fifo_mul_9_32_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_33_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_34_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_35_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_36_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_37_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_38_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_39_ext_size (clk);
            //6� riga
            write_interface #(7,FLUX) wr_fifo_mul_9_40_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_41_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_42_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_43_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_44_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_45_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_46_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_47_ext_size (clk);                        
            //7� riga
            write_interface #(7,FLUX) wr_fifo_mul_9_48_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_49_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_50_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_51_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_52_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_53_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_54_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_55_ext_size (clk);
            //8� riga
            write_interface #(7,FLUX) wr_fifo_mul_9_56_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_57_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_58_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_59_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_60_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_61_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_62_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_9_63_ext_size (clk);
            
            //REMOVE H (x1)
            write_interface #(7,FLUX) wr_fifo_remove_h_0_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_h_1_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_h_2_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_h_3_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_h_4_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_h_5_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_h_6_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_h_7_ext_size (clk);
			
            
            //MUL18 (x64)
            
            //1� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_0_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_1_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_2_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_3_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_4_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_5_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_6_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_7_ext_size (clk);
            //2� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_8_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_9_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_10_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_11_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_12_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_13_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_14_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_15_ext_size (clk);            
            //3� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_16_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_17_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_18_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_19_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_20_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_21_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_22_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_23_ext_size (clk);
            //4� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_24_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_25_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_26_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_27_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_28_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_29_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_30_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_31_ext_size (clk);
            //5� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_32_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_33_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_34_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_35_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_36_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_37_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_38_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_39_ext_size (clk);
            //6� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_40_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_41_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_42_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_43_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_44_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_45_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_46_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_47_ext_size (clk);                        
            //7� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_48_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_49_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_50_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_51_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_52_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_53_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_54_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_55_ext_size (clk);
            //8� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_56_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_57_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_58_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_59_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_60_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_61_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_62_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_63_ext_size (clk);
            
            //REMOVE V (x1)
            write_interface #(7,FLUX) wr_fifo_remove_v_0_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_1_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_2_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_3_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_4_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_5_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_6_ext_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_7_ext_size (clk);
            
            //LINE BUFFER (x7)
            write_interface #(7,FLUX) wr_fifo_line_buffer_0_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_1_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_2_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_3_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_4_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_5_ext_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_6_ext_size (clk);            
                                    
            //DERIVE REAL SIZE (x1)
            write_interface #(7,FLUX) wr_fifo_derive_real_size_ext_size (clk);
                        
        // - FULL            
            assign write_port_ext_size.full =
            
            //MUL9 (x64)
            //1� riga
             wr_fifo_mul_9_0_ext_size.full |
             wr_fifo_mul_9_1_ext_size.full |
             wr_fifo_mul_9_2_ext_size.full |
             wr_fifo_mul_9_3_ext_size.full |
             wr_fifo_mul_9_4_ext_size.full |
             wr_fifo_mul_9_5_ext_size.full |
             wr_fifo_mul_9_6_ext_size.full |
             wr_fifo_mul_9_7_ext_size.full |
            //2� riga
             wr_fifo_mul_9_8_ext_size.full |
             wr_fifo_mul_9_9_ext_size.full |
             wr_fifo_mul_9_10_ext_size.full |
             wr_fifo_mul_9_11_ext_size.full |
             wr_fifo_mul_9_12_ext_size.full |
             wr_fifo_mul_9_13_ext_size.full |
             wr_fifo_mul_9_14_ext_size.full |
             wr_fifo_mul_9_15_ext_size.full |            
            //3� riga
             wr_fifo_mul_9_16_ext_size.full |
             wr_fifo_mul_9_17_ext_size.full |
             wr_fifo_mul_9_18_ext_size.full |
             wr_fifo_mul_9_19_ext_size.full |
             wr_fifo_mul_9_20_ext_size.full |
             wr_fifo_mul_9_21_ext_size.full |
             wr_fifo_mul_9_22_ext_size.full |
             wr_fifo_mul_9_23_ext_size.full |
            //4� riga
             wr_fifo_mul_9_24_ext_size.full |
             wr_fifo_mul_9_25_ext_size.full |
             wr_fifo_mul_9_26_ext_size.full |
             wr_fifo_mul_9_27_ext_size.full |
             wr_fifo_mul_9_28_ext_size.full |
             wr_fifo_mul_9_29_ext_size.full |
             wr_fifo_mul_9_30_ext_size.full |
             wr_fifo_mul_9_31_ext_size.full |
            //5� riga
             wr_fifo_mul_9_32_ext_size.full |
             wr_fifo_mul_9_33_ext_size.full |
             wr_fifo_mul_9_34_ext_size.full |
             wr_fifo_mul_9_35_ext_size.full |
             wr_fifo_mul_9_36_ext_size.full |
             wr_fifo_mul_9_37_ext_size.full |
             wr_fifo_mul_9_38_ext_size.full |
             wr_fifo_mul_9_39_ext_size.full |
            //6� riga
             wr_fifo_mul_9_40_ext_size.full |
             wr_fifo_mul_9_41_ext_size.full |
             wr_fifo_mul_9_42_ext_size.full |
             wr_fifo_mul_9_43_ext_size.full |
             wr_fifo_mul_9_44_ext_size.full |
             wr_fifo_mul_9_45_ext_size.full |
             wr_fifo_mul_9_46_ext_size.full |
             wr_fifo_mul_9_47_ext_size.full |                        
            //7� riga
             wr_fifo_mul_9_48_ext_size.full |
             wr_fifo_mul_9_49_ext_size.full |
             wr_fifo_mul_9_50_ext_size.full |
             wr_fifo_mul_9_51_ext_size.full |
             wr_fifo_mul_9_52_ext_size.full |
             wr_fifo_mul_9_53_ext_size.full |
             wr_fifo_mul_9_54_ext_size.full |
             wr_fifo_mul_9_55_ext_size.full |
            //8� riga
             wr_fifo_mul_9_56_ext_size.full |
             wr_fifo_mul_9_57_ext_size.full |
             wr_fifo_mul_9_58_ext_size.full |
             wr_fifo_mul_9_59_ext_size.full |
             wr_fifo_mul_9_60_ext_size.full |
             wr_fifo_mul_9_61_ext_size.full |
             wr_fifo_mul_9_62_ext_size.full |
             wr_fifo_mul_9_63_ext_size.full |
            
            //REMOVE H (x1)
            wr_fifo_remove_h_0_ext_size.full |
			wr_fifo_remove_h_1_ext_size.full |
			wr_fifo_remove_h_2_ext_size.full |
			wr_fifo_remove_h_3_ext_size.full |
			wr_fifo_remove_h_4_ext_size.full |
			wr_fifo_remove_h_5_ext_size.full |
			wr_fifo_remove_h_6_ext_size.full |
			wr_fifo_remove_h_7_ext_size.full |
            
            //MUL18 (x64)
            //1� riga
             wr_fifo_mul_18_0_ext_size.full |
             wr_fifo_mul_18_1_ext_size.full |
             wr_fifo_mul_18_2_ext_size.full |
             wr_fifo_mul_18_3_ext_size.full |
             wr_fifo_mul_18_4_ext_size.full |
             wr_fifo_mul_18_5_ext_size.full |
             wr_fifo_mul_18_6_ext_size.full |
             wr_fifo_mul_18_7_ext_size.full |
            //2� riga
             wr_fifo_mul_18_8_ext_size.full |
             wr_fifo_mul_18_9_ext_size.full |
             wr_fifo_mul_18_10_ext_size.full |
             wr_fifo_mul_18_11_ext_size.full |
             wr_fifo_mul_18_12_ext_size.full |
             wr_fifo_mul_18_13_ext_size.full |
             wr_fifo_mul_18_14_ext_size.full |
             wr_fifo_mul_18_15_ext_size.full |            
            //3� riga
             wr_fifo_mul_18_16_ext_size.full |
             wr_fifo_mul_18_17_ext_size.full |
             wr_fifo_mul_18_18_ext_size.full |
             wr_fifo_mul_18_19_ext_size.full |
             wr_fifo_mul_18_20_ext_size.full |
             wr_fifo_mul_18_21_ext_size.full |
             wr_fifo_mul_18_22_ext_size.full |
             wr_fifo_mul_18_23_ext_size.full |
            //4� riga
             wr_fifo_mul_18_24_ext_size.full |
             wr_fifo_mul_18_25_ext_size.full |
             wr_fifo_mul_18_26_ext_size.full |
             wr_fifo_mul_18_27_ext_size.full |
             wr_fifo_mul_18_28_ext_size.full |
             wr_fifo_mul_18_29_ext_size.full |
             wr_fifo_mul_18_30_ext_size.full |
             wr_fifo_mul_18_31_ext_size.full |
            //5� riga
             wr_fifo_mul_18_32_ext_size.full |
             wr_fifo_mul_18_33_ext_size.full |
             wr_fifo_mul_18_34_ext_size.full |
             wr_fifo_mul_18_35_ext_size.full |
             wr_fifo_mul_18_36_ext_size.full |
             wr_fifo_mul_18_37_ext_size.full |
             wr_fifo_mul_18_38_ext_size.full |
             wr_fifo_mul_18_39_ext_size.full |
            //6� riga
             wr_fifo_mul_18_40_ext_size.full |
             wr_fifo_mul_18_41_ext_size.full |
             wr_fifo_mul_18_42_ext_size.full |
             wr_fifo_mul_18_43_ext_size.full |
             wr_fifo_mul_18_44_ext_size.full |
             wr_fifo_mul_18_45_ext_size.full |
             wr_fifo_mul_18_46_ext_size.full |
             wr_fifo_mul_18_47_ext_size.full |                        
            //7� riga
             wr_fifo_mul_18_48_ext_size.full |
             wr_fifo_mul_18_49_ext_size.full |
             wr_fifo_mul_18_50_ext_size.full |
             wr_fifo_mul_18_51_ext_size.full |
             wr_fifo_mul_18_52_ext_size.full |
             wr_fifo_mul_18_53_ext_size.full |
             wr_fifo_mul_18_54_ext_size.full |
             wr_fifo_mul_18_55_ext_size.full |
            //8� riga
             wr_fifo_mul_18_56_ext_size.full |
             wr_fifo_mul_18_57_ext_size.full |
             wr_fifo_mul_18_58_ext_size.full |
             wr_fifo_mul_18_59_ext_size.full |
             wr_fifo_mul_18_60_ext_size.full |
             wr_fifo_mul_18_61_ext_size.full |
             wr_fifo_mul_18_62_ext_size.full |
             wr_fifo_mul_18_63_ext_size.full |
            
            //REMOVE V (x1)
            wr_fifo_remove_v_0_ext_size.full |
			wr_fifo_remove_v_1_ext_size.full |
			wr_fifo_remove_v_2_ext_size.full |
			wr_fifo_remove_v_3_ext_size.full |
			wr_fifo_remove_v_4_ext_size.full |
			wr_fifo_remove_v_5_ext_size.full |
			wr_fifo_remove_v_6_ext_size.full |
			wr_fifo_remove_v_7_ext_size.full |
            
            //LINE BUFFER (x7)
            wr_fifo_line_buffer_0_ext_size.full |
            wr_fifo_line_buffer_1_ext_size.full |
            wr_fifo_line_buffer_2_ext_size.full |
            wr_fifo_line_buffer_3_ext_size.full |
            wr_fifo_line_buffer_4_ext_size.full |
            wr_fifo_line_buffer_5_ext_size.full |
            wr_fifo_line_buffer_6_ext_size.full |            
                                    
            //DERIVE REAL SIZE (x1)
            wr_fifo_derive_real_size_ext_size.full ;             
                        
        // - WRITE
            
            //MUL9 (x64) 
            //1� riga
             assign wr_fifo_mul_9_0_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_1_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_2_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_3_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_4_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_5_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_6_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_7_ext_size.write = write_port_ext_size.write;
            //2� riga
             assign wr_fifo_mul_9_8_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_9_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_10_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_11_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_12_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_13_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_14_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_15_ext_size.write = write_port_ext_size.write;            
            //3� riga
             assign wr_fifo_mul_9_16_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_17_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_18_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_19_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_20_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_21_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_22_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_23_ext_size.write = write_port_ext_size.write;
            //4� riga
             assign wr_fifo_mul_9_24_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_25_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_26_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_27_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_28_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_29_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_30_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_31_ext_size.write = write_port_ext_size.write;
            //5� riga
             assign wr_fifo_mul_9_32_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_33_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_34_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_35_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_36_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_37_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_38_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_39_ext_size.write = write_port_ext_size.write;
            //6� riga
             assign wr_fifo_mul_9_40_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_41_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_42_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_43_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_44_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_45_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_46_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_47_ext_size.write = write_port_ext_size.write;
            //7� riga
             assign wr_fifo_mul_9_48_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_49_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_50_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_51_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_52_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_53_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_54_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_55_ext_size.write = write_port_ext_size.write;
            //8� riga
             assign wr_fifo_mul_9_56_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_57_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_58_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_59_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_60_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_61_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_62_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_9_63_ext_size.write = write_port_ext_size.write;
            
            //REMOVE H (x1)
            assign wr_fifo_remove_h_0_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_h_1_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_h_2_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_h_3_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_h_4_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_h_5_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_h_6_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_h_7_ext_size.write = write_port_ext_size.write;

			
            
            //MUL18 (x64)
            //1� riga
             assign wr_fifo_mul_18_0_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_1_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_2_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_3_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_4_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_5_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_6_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_7_ext_size.write = write_port_ext_size.write;
            //2� riga
             assign wr_fifo_mul_18_8_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_9_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_10_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_11_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_12_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_13_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_14_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_15_ext_size.write = write_port_ext_size.write;            
            //3� riga
             assign wr_fifo_mul_18_16_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_17_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_18_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_19_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_20_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_21_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_22_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_23_ext_size.write = write_port_ext_size.write;
            //4� riga
             assign wr_fifo_mul_18_24_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_25_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_26_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_27_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_28_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_29_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_30_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_31_ext_size.write = write_port_ext_size.write;
            //5� riga
             assign wr_fifo_mul_18_32_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_33_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_34_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_35_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_36_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_37_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_38_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_39_ext_size.write = write_port_ext_size.write;
            //6� riga
             assign wr_fifo_mul_18_40_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_41_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_42_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_43_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_44_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_45_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_46_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_47_ext_size.write = write_port_ext_size.write;
            //7� riga
             assign wr_fifo_mul_18_48_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_49_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_50_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_51_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_52_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_53_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_54_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_55_ext_size.write = write_port_ext_size.write;
            //8� riga
             assign wr_fifo_mul_18_56_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_57_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_58_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_59_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_60_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_61_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_62_ext_size.write = write_port_ext_size.write;
             assign wr_fifo_mul_18_63_ext_size.write = write_port_ext_size.write;
            
            //REMOVE V (x1)
            assign wr_fifo_remove_v_0_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_v_1_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_v_2_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_v_3_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_v_4_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_v_5_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_v_6_ext_size.write = write_port_ext_size.write;
			assign wr_fifo_remove_v_7_ext_size.write = write_port_ext_size.write;
            
            //LINE BUFFER (x7)
            assign wr_fifo_line_buffer_0_ext_size.write = write_port_ext_size.write;
            assign wr_fifo_line_buffer_1_ext_size.write = write_port_ext_size.write;
            assign wr_fifo_line_buffer_2_ext_size.write = write_port_ext_size.write;
            assign wr_fifo_line_buffer_3_ext_size.write = write_port_ext_size.write;
            assign wr_fifo_line_buffer_4_ext_size.write = write_port_ext_size.write;
            assign wr_fifo_line_buffer_5_ext_size.write = write_port_ext_size.write;
            assign wr_fifo_line_buffer_6_ext_size.write = write_port_ext_size.write;            
                                    
            //DERIVE REAL SIZE (x1)
            assign wr_fifo_derive_real_size_ext_size.write = write_port_ext_size.write; 
                        
        // - DATA
            
            //MUL9 (x64) 
            //1� riga
             assign wr_fifo_mul_9_0_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_1_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_2_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_3_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_4_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_5_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_6_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_7_ext_size.din = write_port_ext_size.din;
            //2� riga
             assign wr_fifo_mul_9_8_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_9_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_10_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_11_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_12_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_13_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_14_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_15_ext_size.din = write_port_ext_size.din;            
            //3� riga
             assign wr_fifo_mul_9_16_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_17_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_18_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_19_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_20_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_21_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_22_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_23_ext_size.din = write_port_ext_size.din;
            //4� riga
             assign wr_fifo_mul_9_24_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_25_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_26_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_27_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_28_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_29_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_30_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_31_ext_size.din = write_port_ext_size.din;
            //5� riga
             assign wr_fifo_mul_9_32_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_33_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_34_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_35_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_36_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_37_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_38_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_39_ext_size.din = write_port_ext_size.din;
            //6� riga
             assign wr_fifo_mul_9_40_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_41_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_42_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_43_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_44_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_45_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_46_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_47_ext_size.din = write_port_ext_size.din;
            //7� riga
             assign wr_fifo_mul_9_48_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_49_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_50_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_51_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_52_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_53_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_54_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_55_ext_size.din = write_port_ext_size.din;
            //8� riga
             assign wr_fifo_mul_9_56_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_57_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_58_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_59_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_60_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_61_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_62_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_9_63_ext_size.din = write_port_ext_size.din;
            
            //REMOVE H (x1)
            assign wr_fifo_remove_h_0_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_h_1_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_h_2_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_h_3_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_h_4_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_h_5_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_h_6_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_h_7_ext_size.din = write_port_ext_size.din;
            
            //MUL18 (x64)
            //1� riga
             assign wr_fifo_mul_18_0_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_1_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_2_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_3_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_4_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_5_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_6_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_7_ext_size.din = write_port_ext_size.din;
            //2� riga
             assign wr_fifo_mul_18_8_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_9_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_10_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_11_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_12_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_13_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_14_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_15_ext_size.din = write_port_ext_size.din;            
            //3� riga
             assign wr_fifo_mul_18_16_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_17_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_18_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_19_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_20_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_21_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_22_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_23_ext_size.din = write_port_ext_size.din;
            //4� riga
             assign wr_fifo_mul_18_24_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_25_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_26_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_27_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_28_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_29_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_30_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_31_ext_size.din = write_port_ext_size.din;
            //5� riga
             assign wr_fifo_mul_18_32_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_33_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_34_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_35_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_36_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_37_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_38_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_39_ext_size.din = write_port_ext_size.din;
            //6� riga
             assign wr_fifo_mul_18_40_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_41_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_42_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_43_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_44_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_45_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_46_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_47_ext_size.din = write_port_ext_size.din;
            //7� riga
             assign wr_fifo_mul_18_48_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_49_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_50_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_51_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_52_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_53_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_54_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_55_ext_size.din = write_port_ext_size.din;
            //8� riga
             assign wr_fifo_mul_18_56_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_57_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_58_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_59_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_60_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_61_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_62_ext_size.din = write_port_ext_size.din;
             assign wr_fifo_mul_18_63_ext_size.din = write_port_ext_size.din;
            
            //REMOVE V (x1)
            assign wr_fifo_remove_v_0_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_v_1_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_v_2_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_v_3_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_v_4_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_v_5_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_v_6_ext_size.din = write_port_ext_size.din;
			assign wr_fifo_remove_v_7_ext_size.din = write_port_ext_size.din;
            
            //LINE BUFFER (x7)
            assign wr_fifo_line_buffer_0_ext_size.din = write_port_ext_size.din;
            assign wr_fifo_line_buffer_1_ext_size.din = write_port_ext_size.din;
            assign wr_fifo_line_buffer_2_ext_size.din = write_port_ext_size.din;
            assign wr_fifo_line_buffer_3_ext_size.din = write_port_ext_size.din;
            assign wr_fifo_line_buffer_4_ext_size.din = write_port_ext_size.din;
            assign wr_fifo_line_buffer_5_ext_size.din = write_port_ext_size.din;
            assign wr_fifo_line_buffer_6_ext_size.din = write_port_ext_size.din;            
                                    
            //DERIVE REAL SIZE (x1)
            assign wr_fifo_derive_real_size_ext_size.din = write_port_ext_size.din;

    //FORK LINE_BUFFER_0 / LINE_BUFFER_1 / LINE_BUFFER_2 / LINE_BUFFER_3 / LINE_BUFFER_4 ...
    //... / LINE_BUFFER_5 / LINE_BUFFER_6  / REMOVE_V / MUL_18_0 / MUL_18_1 / MUL_18_2 ... 
    //... / MUL_18_3 / MUL_18_4 / MUL_18_5 / MUL_18_6 / MUL_18_7...
    //... ON DERIVE_REAL_SIZE 

        // - INTERFACES
            
            //MUL18 (x64)
            //1� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_0_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_1_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_2_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_3_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_4_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_5_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_6_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_7_real_size (clk);
            //2� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_8_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_9_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_10_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_11_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_12_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_13_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_14_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_15_real_size (clk);            
            //3� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_16_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_17_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_18_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_19_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_20_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_21_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_22_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_23_real_size (clk);
            //4� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_24_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_25_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_26_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_27_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_28_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_29_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_30_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_31_real_size (clk);
            //5� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_32_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_33_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_34_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_35_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_36_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_37_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_38_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_39_real_size (clk);
            //6� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_40_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_41_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_42_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_43_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_44_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_45_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_46_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_47_real_size (clk);                        
            //7� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_48_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_49_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_50_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_51_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_52_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_53_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_54_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_55_real_size (clk);
            //8� riga
            write_interface #(7,FLUX) wr_fifo_mul_18_56_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_57_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_58_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_59_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_60_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_61_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_62_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_mul_18_63_real_size (clk);
            
            //REMOVE V (x1)
            write_interface #(7,FLUX) wr_fifo_remove_v_0_real_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_1_real_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_2_real_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_3_real_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_4_real_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_5_real_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_6_real_size (clk);
			write_interface #(7,FLUX) wr_fifo_remove_v_7_real_size (clk);
            
            //LINE BUFFER (x7)
            write_interface #(7,FLUX) wr_fifo_line_buffer_0_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_1_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_2_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_3_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_4_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_5_real_size (clk);
            write_interface #(7,FLUX) wr_fifo_line_buffer_6_real_size (clk);            
                                                          
        // - FULL            
            assign wr_derive_real_size_real_size.full =
            
            //MUL18 (x64)
            //1� riga
             wr_fifo_mul_18_0_real_size.full |
             wr_fifo_mul_18_1_real_size.full |
             wr_fifo_mul_18_2_real_size.full |
             wr_fifo_mul_18_3_real_size.full |
             wr_fifo_mul_18_4_real_size.full |
             wr_fifo_mul_18_5_real_size.full |
             wr_fifo_mul_18_6_real_size.full |
             wr_fifo_mul_18_7_real_size.full |
            //2� riga
             wr_fifo_mul_18_8_real_size.full |
             wr_fifo_mul_18_9_real_size.full |
             wr_fifo_mul_18_10_real_size.full |
             wr_fifo_mul_18_11_real_size.full |
             wr_fifo_mul_18_12_real_size.full |
             wr_fifo_mul_18_13_real_size.full |
             wr_fifo_mul_18_14_real_size.full |
             wr_fifo_mul_18_15_real_size.full |            
            //3� riga
             wr_fifo_mul_18_16_real_size.full |
             wr_fifo_mul_18_17_real_size.full |
             wr_fifo_mul_18_18_real_size.full |
             wr_fifo_mul_18_19_real_size.full |
             wr_fifo_mul_18_20_real_size.full |
             wr_fifo_mul_18_21_real_size.full |
             wr_fifo_mul_18_22_real_size.full |
             wr_fifo_mul_18_23_real_size.full |
            //4� riga
             wr_fifo_mul_18_24_real_size.full |
             wr_fifo_mul_18_25_real_size.full |
             wr_fifo_mul_18_26_real_size.full |
             wr_fifo_mul_18_27_real_size.full |
             wr_fifo_mul_18_28_real_size.full |
             wr_fifo_mul_18_29_real_size.full |
             wr_fifo_mul_18_30_real_size.full |
             wr_fifo_mul_18_31_real_size.full |
            //5� riga
             wr_fifo_mul_18_32_real_size.full |
             wr_fifo_mul_18_33_real_size.full |
             wr_fifo_mul_18_34_real_size.full |
             wr_fifo_mul_18_35_real_size.full |
             wr_fifo_mul_18_36_real_size.full |
             wr_fifo_mul_18_37_real_size.full |
             wr_fifo_mul_18_38_real_size.full |
             wr_fifo_mul_18_39_real_size.full |
            //6� riga
             wr_fifo_mul_18_40_real_size.full |
             wr_fifo_mul_18_41_real_size.full |
             wr_fifo_mul_18_42_real_size.full |
             wr_fifo_mul_18_43_real_size.full |
             wr_fifo_mul_18_44_real_size.full |
             wr_fifo_mul_18_45_real_size.full |
             wr_fifo_mul_18_46_real_size.full |
             wr_fifo_mul_18_47_real_size.full |                        
            //7� riga
             wr_fifo_mul_18_48_real_size.full |
             wr_fifo_mul_18_49_real_size.full |
             wr_fifo_mul_18_50_real_size.full |
             wr_fifo_mul_18_51_real_size.full |
             wr_fifo_mul_18_52_real_size.full |
             wr_fifo_mul_18_53_real_size.full |
             wr_fifo_mul_18_54_real_size.full |
             wr_fifo_mul_18_55_real_size.full |
            //8� riga
             wr_fifo_mul_18_56_real_size.full |
             wr_fifo_mul_18_57_real_size.full |
             wr_fifo_mul_18_58_real_size.full |
             wr_fifo_mul_18_59_real_size.full |
             wr_fifo_mul_18_60_real_size.full |
             wr_fifo_mul_18_61_real_size.full |
             wr_fifo_mul_18_62_real_size.full |
             wr_fifo_mul_18_63_real_size.full |
            
            //REMOVE V (x1)
            wr_fifo_remove_v_0_real_size.full |
			wr_fifo_remove_v_1_real_size.full |
			wr_fifo_remove_v_2_real_size.full |
			wr_fifo_remove_v_3_real_size.full |
			wr_fifo_remove_v_4_real_size.full |
			wr_fifo_remove_v_5_real_size.full |
			wr_fifo_remove_v_6_real_size.full |
			wr_fifo_remove_v_7_real_size.full |
            
            //LINE BUFFER (x7)
            wr_fifo_line_buffer_0_real_size.full |
            wr_fifo_line_buffer_1_real_size.full |
            wr_fifo_line_buffer_2_real_size.full |
            wr_fifo_line_buffer_3_real_size.full |
            wr_fifo_line_buffer_4_real_size.full |
            wr_fifo_line_buffer_5_real_size.full |
            wr_fifo_line_buffer_6_real_size.full ;            
                                                              
        // - WRITE
                        
            //MUL18 (x8)
            //1� riga
             assign wr_fifo_mul_18_0_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_1_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_2_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_3_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_4_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_5_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_6_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_7_real_size.write = wr_derive_real_size_real_size.write;
            //2� riga
             assign wr_fifo_mul_18_8_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_9_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_10_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_11_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_12_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_13_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_14_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_15_real_size.write = wr_derive_real_size_real_size.write;            
            //3� riga
             assign wr_fifo_mul_18_16_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_17_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_18_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_19_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_20_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_21_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_22_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_23_real_size.write = wr_derive_real_size_real_size.write;
            //4� riga
             assign wr_fifo_mul_18_24_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_25_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_26_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_27_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_28_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_29_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_30_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_31_real_size.write = wr_derive_real_size_real_size.write;
            //5� riga
             assign wr_fifo_mul_18_32_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_33_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_34_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_35_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_36_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_37_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_38_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_39_real_size.write = wr_derive_real_size_real_size.write;
            //6� riga
             assign wr_fifo_mul_18_40_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_41_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_42_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_43_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_44_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_45_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_46_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_47_real_size.write = wr_derive_real_size_real_size.write;
            //7� riga
             assign wr_fifo_mul_18_48_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_49_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_50_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_51_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_52_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_53_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_54_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_55_real_size.write = wr_derive_real_size_real_size.write;
            //8� riga
             assign wr_fifo_mul_18_56_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_57_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_58_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_59_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_60_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_61_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_62_real_size.write = wr_derive_real_size_real_size.write;
             assign wr_fifo_mul_18_63_real_size.write = wr_derive_real_size_real_size.write;
            
            //REMOVE V (x1)
            assign wr_fifo_remove_v_0_real_size.write = wr_derive_real_size_real_size.write;
			assign wr_fifo_remove_v_1_real_size.write = wr_derive_real_size_real_size.write;
			assign wr_fifo_remove_v_2_real_size.write = wr_derive_real_size_real_size.write;
			assign wr_fifo_remove_v_3_real_size.write = wr_derive_real_size_real_size.write;
			assign wr_fifo_remove_v_4_real_size.write = wr_derive_real_size_real_size.write;
			assign wr_fifo_remove_v_5_real_size.write = wr_derive_real_size_real_size.write;
			assign wr_fifo_remove_v_6_real_size.write = wr_derive_real_size_real_size.write;
			assign wr_fifo_remove_v_7_real_size.write = wr_derive_real_size_real_size.write;
            
            //LINE BUFFER (x7)
            assign wr_fifo_line_buffer_0_real_size.write = wr_derive_real_size_real_size.write;
            assign wr_fifo_line_buffer_1_real_size.write = wr_derive_real_size_real_size.write;
            assign wr_fifo_line_buffer_2_real_size.write = wr_derive_real_size_real_size.write;
            assign wr_fifo_line_buffer_3_real_size.write = wr_derive_real_size_real_size.write;
            assign wr_fifo_line_buffer_4_real_size.write = wr_derive_real_size_real_size.write;
            assign wr_fifo_line_buffer_5_real_size.write = wr_derive_real_size_real_size.write;
            assign wr_fifo_line_buffer_6_real_size.write = wr_derive_real_size_real_size.write;            
                    
        // - DATA
                                
            //MUL18 (x8)
            //1� riga
             assign wr_fifo_mul_18_0_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_1_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_2_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_3_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_4_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_5_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_6_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_7_real_size.din = wr_derive_real_size_real_size.din;
            //2� riga
             assign wr_fifo_mul_18_8_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_9_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_10_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_11_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_12_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_13_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_14_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_15_real_size.din = wr_derive_real_size_real_size.din;            
            //3� riga
             assign wr_fifo_mul_18_16_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_17_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_18_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_19_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_20_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_21_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_22_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_23_real_size.din = wr_derive_real_size_real_size.din;
            //4� riga
             assign wr_fifo_mul_18_24_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_25_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_26_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_27_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_28_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_29_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_30_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_31_real_size.din = wr_derive_real_size_real_size.din;
            //5� riga
             assign wr_fifo_mul_18_32_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_33_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_34_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_35_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_36_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_37_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_38_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_39_real_size.din = wr_derive_real_size_real_size.din;
            //6� riga
             assign wr_fifo_mul_18_40_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_41_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_42_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_43_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_44_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_45_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_46_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_47_real_size.din = wr_derive_real_size_real_size.din;
            //7� riga
             assign wr_fifo_mul_18_48_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_49_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_50_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_51_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_52_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_53_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_54_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_55_real_size.din = wr_derive_real_size_real_size.din;
            //8� riga
             assign wr_fifo_mul_18_56_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_57_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_58_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_59_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_60_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_61_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_62_real_size.din = wr_derive_real_size_real_size.din;
             assign wr_fifo_mul_18_63_real_size.din = wr_derive_real_size_real_size.din;
            
            //REMOVE V (x1)
            assign wr_fifo_remove_v_0_real_size.din = wr_derive_real_size_real_size.din;
			assign wr_fifo_remove_v_1_real_size.din = wr_derive_real_size_real_size.din;
			assign wr_fifo_remove_v_2_real_size.din = wr_derive_real_size_real_size.din;
			assign wr_fifo_remove_v_3_real_size.din = wr_derive_real_size_real_size.din;
			assign wr_fifo_remove_v_4_real_size.din = wr_derive_real_size_real_size.din;
			assign wr_fifo_remove_v_5_real_size.din = wr_derive_real_size_real_size.din;
			assign wr_fifo_remove_v_6_real_size.din = wr_derive_real_size_real_size.din;
			assign wr_fifo_remove_v_7_real_size.din = wr_derive_real_size_real_size.din;
            
            //LINE BUFFER (x7)
            assign wr_fifo_line_buffer_0_real_size.din = wr_derive_real_size_real_size.din;
            assign wr_fifo_line_buffer_1_real_size.din = wr_derive_real_size_real_size.din;
            assign wr_fifo_line_buffer_2_real_size.din = wr_derive_real_size_real_size.din;
            assign wr_fifo_line_buffer_3_real_size.din = wr_derive_real_size_real_size.din;
            assign wr_fifo_line_buffer_4_real_size.din = wr_derive_real_size_real_size.din;
            assign wr_fifo_line_buffer_5_real_size.din = wr_derive_real_size_real_size.din;
            assign wr_fifo_line_buffer_6_real_size.din = wr_derive_real_size_real_size.din; 


    //FORK INPUT 0 TO MUL_9_0 & MUL_9_15 & MUL_9_22 & MUL_9_29 & MUL_9_36 & MUL_9_43 & MUL_9_50 & MUL_9_57

        // - INTERFACES   		
        write_interface #(8,FLUX) wr_fifo_mul_9_0_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_15_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_22_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_29_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_36_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_43_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_50_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_57_opA(clk); 
               
        // - FULL
        assign write_port_in_port_0.full = wr_fifo_mul_9_0_opA.full 
        | wr_fifo_mul_9_15_opA.full | wr_fifo_mul_9_22_opA.full | wr_fifo_mul_9_29_opA.full | wr_fifo_mul_9_36_opA.full
        | wr_fifo_mul_9_43_opA.full | wr_fifo_mul_9_50_opA.full | wr_fifo_mul_9_57_opA.full;
        
        // - WRITE
        assign wr_fifo_mul_9_0_opA.write = write_port_in_port_0.write;
        assign wr_fifo_mul_9_15_opA.write = write_port_in_port_0.write;
        assign wr_fifo_mul_9_22_opA.write = write_port_in_port_0.write;
        assign wr_fifo_mul_9_29_opA.write = write_port_in_port_0.write;
        assign wr_fifo_mul_9_36_opA.write = write_port_in_port_0.write;
        assign wr_fifo_mul_9_43_opA.write = write_port_in_port_0.write;
        assign wr_fifo_mul_9_50_opA.write = write_port_in_port_0.write;
        assign wr_fifo_mul_9_57_opA.write = write_port_in_port_0.write;
        
        // - DATA
        assign wr_fifo_mul_9_0_opA.din = write_port_in_port_0.din;
        assign wr_fifo_mul_9_15_opA.din = write_port_in_port_0.din;
        assign wr_fifo_mul_9_22_opA.din = write_port_in_port_0.din;
        assign wr_fifo_mul_9_29_opA.din = write_port_in_port_0.din;
        assign wr_fifo_mul_9_36_opA.din = write_port_in_port_0.din;
        assign wr_fifo_mul_9_43_opA.din = write_port_in_port_0.din;
        assign wr_fifo_mul_9_50_opA.din = write_port_in_port_0.din;
        assign wr_fifo_mul_9_57_opA.din = write_port_in_port_0.din;
    
    //FORK INPUT 1 TO DELAY_0 & MUL_9_1 & MUL_9_23 & MUL_9_30 & MUL_9_37 & MUL_9_44 & MUL_9_51 & MUL_9_58 

        // - INTERFACES   		
        write_interface #(8,FLUX) wr_fifo_delay_0_in_pel(clk);    		
        write_interface #(8,FLUX) wr_fifo_mul_9_1_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_23_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_30_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_37_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_44_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_51_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_58_opA(clk); 
               
        // - FULL
        assign write_port_in_port_1.full = wr_fifo_delay_0_in_pel.full | wr_fifo_mul_9_1_opA.full 
        | wr_fifo_mul_9_23_opA.full | wr_fifo_mul_9_30_opA.full | wr_fifo_mul_9_37_opA.full
        | wr_fifo_mul_9_44_opA.full | wr_fifo_mul_9_51_opA.full | wr_fifo_mul_9_58_opA.full;
        
        // - WRITE
        assign wr_fifo_delay_0_in_pel.write = write_port_in_port_1.write;
        assign wr_fifo_mul_9_1_opA.write = write_port_in_port_1.write;
        assign wr_fifo_mul_9_23_opA.write = write_port_in_port_1.write;
        assign wr_fifo_mul_9_30_opA.write = write_port_in_port_1.write;
        assign wr_fifo_mul_9_37_opA.write = write_port_in_port_1.write;
        assign wr_fifo_mul_9_44_opA.write = write_port_in_port_1.write;
        assign wr_fifo_mul_9_51_opA.write = write_port_in_port_1.write;
        assign wr_fifo_mul_9_58_opA.write = write_port_in_port_1.write;
        
        // - DATA
        assign wr_fifo_delay_0_in_pel.din = write_port_in_port_1.din;
        assign wr_fifo_mul_9_1_opA.din = write_port_in_port_1.din;
        assign wr_fifo_mul_9_23_opA.din = write_port_in_port_1.din;
        assign wr_fifo_mul_9_30_opA.din = write_port_in_port_1.din;
        assign wr_fifo_mul_9_37_opA.din = write_port_in_port_1.din;
        assign wr_fifo_mul_9_44_opA.din = write_port_in_port_1.din;
        assign wr_fifo_mul_9_51_opA.din = write_port_in_port_1.din;
        assign wr_fifo_mul_9_58_opA.din = write_port_in_port_1.din;


	//FORK INPUT 2 TO DELAY_1 & MUL_9_2 & MUL_9_31 & MUL_9_38 & MUL_9_45 & MUL_9_52 & MUL_9_59
	
        // - INTERFACES   		
        write_interface #(8,FLUX) wr_fifo_delay_1_in_pel(clk);    		
        write_interface #(8,FLUX) wr_fifo_mul_9_2_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_31_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_38_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_45_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_52_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_59_opA(clk); 
               
        // - FULL
        assign write_port_in_port_2.full = wr_fifo_delay_1_in_pel.full | wr_fifo_mul_9_2_opA.full 
        | wr_fifo_mul_9_31_opA.full | wr_fifo_mul_9_38_opA.full
        | wr_fifo_mul_9_45_opA.full | wr_fifo_mul_9_52_opA.full | wr_fifo_mul_9_59_opA.full;
        
        // - WRITE
        assign wr_fifo_delay_1_in_pel.write = write_port_in_port_2.write;
        assign wr_fifo_mul_9_2_opA.write = write_port_in_port_2.write;
        assign wr_fifo_mul_9_31_opA.write = write_port_in_port_2.write;
        assign wr_fifo_mul_9_38_opA.write = write_port_in_port_2.write;
        assign wr_fifo_mul_9_45_opA.write = write_port_in_port_2.write;
        assign wr_fifo_mul_9_52_opA.write = write_port_in_port_2.write;
        assign wr_fifo_mul_9_59_opA.write = write_port_in_port_2.write;
        
        // - DATA
        assign wr_fifo_delay_1_in_pel.din = write_port_in_port_2.din;
        assign wr_fifo_mul_9_2_opA.din = write_port_in_port_2.din;
        assign wr_fifo_mul_9_31_opA.din = write_port_in_port_2.din;
        assign wr_fifo_mul_9_38_opA.din = write_port_in_port_2.din;
        assign wr_fifo_mul_9_45_opA.din = write_port_in_port_2.din;
        assign wr_fifo_mul_9_52_opA.din = write_port_in_port_2.din;
        assign wr_fifo_mul_9_59_opA.din = write_port_in_port_2.din;

    //FORK INPUT 3 TO DELAY_2 & MUL_9_3 & MUL_9_39 & MUL_9_46 & MUL_9_53 & MUL_9_60 

        // - INTERFACES   		
        write_interface #(8,FLUX) wr_fifo_delay_2_in_pel(clk);    		
        write_interface #(8,FLUX) wr_fifo_mul_9_3_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_39_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_46_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_53_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_60_opA(clk); 
               
        // - FULL
        assign write_port_in_port_3.full = wr_fifo_delay_2_in_pel.full | wr_fifo_mul_9_3_opA.full 
        | wr_fifo_mul_9_39_opA.full | wr_fifo_mul_9_46_opA.full | wr_fifo_mul_9_53_opA.full | wr_fifo_mul_9_60_opA.full;
        
        // - WRITE
        assign wr_fifo_delay_2_in_pel.write = write_port_in_port_3.write;
        assign wr_fifo_mul_9_3_opA.write = write_port_in_port_3.write;
        assign wr_fifo_mul_9_39_opA.write = write_port_in_port_3.write;
        assign wr_fifo_mul_9_46_opA.write = write_port_in_port_3.write;
        assign wr_fifo_mul_9_53_opA.write = write_port_in_port_3.write;
        assign wr_fifo_mul_9_60_opA.write = write_port_in_port_3.write;
        
        // - DATA
        assign wr_fifo_delay_2_in_pel.din = write_port_in_port_3.din;
        assign wr_fifo_mul_9_3_opA.din = write_port_in_port_3.din;
        assign wr_fifo_mul_9_39_opA.din = write_port_in_port_3.din;
        assign wr_fifo_mul_9_46_opA.din = write_port_in_port_3.din;
        assign wr_fifo_mul_9_53_opA.din = write_port_in_port_3.din;
        assign wr_fifo_mul_9_60_opA.din = write_port_in_port_3.din;
    
    //FORK INPUT 4 TO DELAY_3 & MUL_9_4 & MUL_9_47 & MUL_9_54 & MUL_9_61
    
        // - INTERFACES   		
        write_interface #(8,FLUX) wr_fifo_delay_3_in_pel(clk);    		
        write_interface #(8,FLUX) wr_fifo_mul_9_4_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_47_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_54_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_61_opA(clk); 
               
        // - FULL
        assign write_port_in_port_4.full = wr_fifo_delay_3_in_pel.full | wr_fifo_mul_9_4_opA.full 
        | wr_fifo_mul_9_47_opA.full | wr_fifo_mul_9_54_opA.full | wr_fifo_mul_9_61_opA.full;
        
        // - WRITE
        assign wr_fifo_delay_3_in_pel.write = write_port_in_port_4.write;
        assign wr_fifo_mul_9_4_opA.write = write_port_in_port_4.write;
        assign wr_fifo_mul_9_47_opA.write = write_port_in_port_4.write;
        assign wr_fifo_mul_9_54_opA.write = write_port_in_port_4.write;
        assign wr_fifo_mul_9_61_opA.write = write_port_in_port_4.write;
        
        // - DATA
        assign wr_fifo_delay_3_in_pel.din = write_port_in_port_4.din;
        assign wr_fifo_mul_9_4_opA.din = write_port_in_port_4.din;
        assign wr_fifo_mul_9_47_opA.din = write_port_in_port_4.din;
        assign wr_fifo_mul_9_54_opA.din = write_port_in_port_4.din;
        assign wr_fifo_mul_9_61_opA.din = write_port_in_port_4.din;
	
    //FORK INPUT 5 TO DELAY_4 & MUL_9_5 & MUL_9_55 & MUL_9_62 

        // - INTERFACES   		
        write_interface #(8,FLUX) wr_fifo_delay_4_in_pel(clk);    		
        write_interface #(8,FLUX) wr_fifo_mul_9_5_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_55_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_62_opA(clk); 
               
        // - FULL
        assign write_port_in_port_5.full = wr_fifo_delay_4_in_pel.full | wr_fifo_mul_9_5_opA.full 
        | wr_fifo_mul_9_55_opA.full | wr_fifo_mul_9_62_opA.full;
        
        // - WRITE
        assign wr_fifo_delay_4_in_pel.write = write_port_in_port_5.write;
        assign wr_fifo_mul_9_5_opA.write = write_port_in_port_5.write;
        assign wr_fifo_mul_9_55_opA.write = write_port_in_port_5.write;
        assign wr_fifo_mul_9_62_opA.write = write_port_in_port_5.write;
        
        // - DATA
        assign wr_fifo_delay_4_in_pel.din = write_port_in_port_5.din;
        assign wr_fifo_mul_9_5_opA.din = write_port_in_port_5.din;
        assign wr_fifo_mul_9_55_opA.din = write_port_in_port_5.din;
        assign wr_fifo_mul_9_62_opA.din = write_port_in_port_5.din;	
    
    //FORK INPUT 6 TO DELAY_5 & MUL_9_6 & MUL_9_63 

        // - INTERFACES   		
        write_interface #(8,FLUX) wr_fifo_delay_5_in_pel(clk);    		
        write_interface #(8,FLUX) wr_fifo_mul_9_6_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_63_opA(clk); 
               
        // - FULL
        assign write_port_in_port_6.full = wr_fifo_delay_5_in_pel.full | wr_fifo_mul_9_6_opA.full 
        | wr_fifo_mul_9_63_opA.full;
        
        // - WRITE
        assign wr_fifo_delay_5_in_pel.write = write_port_in_port_6.write;
        assign wr_fifo_mul_9_6_opA.write = write_port_in_port_6.write;
        assign wr_fifo_mul_9_63_opA.write = write_port_in_port_6.write;
        
        // - DATA
        assign wr_fifo_delay_5_in_pel.din = write_port_in_port_6.din;
        assign wr_fifo_mul_9_6_opA.din = write_port_in_port_6.din;
        assign wr_fifo_mul_9_63_opA.din = write_port_in_port_6.din;	
    
    //FORK INPUT 7 TO DELAY_6 & MUL_9_7 

        // - INTERFACES   		
        write_interface #(8,FLUX) wr_fifo_delay_6_in_pel(clk);    		
        write_interface #(8,FLUX) wr_fifo_mul_9_7_opA(clk);
               
        // - FULL
        assign write_port_in_port_7.full = wr_fifo_delay_6_in_pel.full | wr_fifo_mul_9_7_opA.full;
        
        // - WRITE
        assign wr_fifo_delay_6_in_pel.write = write_port_in_port_7.write;
        assign wr_fifo_mul_9_7_opA.write = write_port_in_port_7.write;
        
        // - DATA
        assign wr_fifo_delay_6_in_pel.din = write_port_in_port_7.din;
        assign wr_fifo_mul_9_7_opA.din = write_port_in_port_7.din;
  
    //FORK DELAY 1 TO MUL_9_9 & MUL_9_16

        // - INTERFACES   		    		
        write_interface #(8,FLUX) wr_fifo_mul_9_9_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_16_opA(clk);
               
        // - FULL
        assign wr_delay_1_out_pel.full = wr_fifo_mul_9_9_opA.full | wr_fifo_mul_9_16_opA.full;
        
        // - WRITE 
        assign wr_fifo_mul_9_9_opA.write = wr_delay_1_out_pel.write;
        assign wr_fifo_mul_9_16_opA.write = wr_delay_1_out_pel.write;
        
        // - DATA
        assign wr_fifo_mul_9_9_opA.din = wr_delay_1_out_pel.din;
        assign wr_fifo_mul_9_16_opA.din = wr_delay_1_out_pel.din;
    
    //FORK DELAY 2 TO MUL_9_10 & MUL_9_17 & MUL_9_24

        // - INTERFACES   		    		
        write_interface #(8,FLUX) wr_fifo_mul_9_10_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_17_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_24_opA(clk);
               
        // - FULL
        assign wr_delay_2_out_pel.full = wr_fifo_mul_9_10_opA.full | wr_fifo_mul_9_17_opA.full | wr_fifo_mul_9_24_opA.full;
        
        // - WRITE 
        assign wr_fifo_mul_9_10_opA.write = wr_delay_2_out_pel.write;
        assign wr_fifo_mul_9_17_opA.write = wr_delay_2_out_pel.write;
        assign wr_fifo_mul_9_24_opA.write = wr_delay_2_out_pel.write;
        
        // - DATA
        assign wr_fifo_mul_9_10_opA.din = wr_delay_2_out_pel.din;
        assign wr_fifo_mul_9_17_opA.din = wr_delay_2_out_pel.din;
        assign wr_fifo_mul_9_24_opA.din = wr_delay_2_out_pel.din;
                    
    //FORK DELAY 3 TO MUL_9_11 & MUL_9_18 & MUL_9_25 & MUL_9_32

        // - INTERFACES   		    		
        write_interface #(8,FLUX) wr_fifo_mul_9_11_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_18_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_25_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_32_opA(clk);
               
        // - FULL
        assign wr_delay_3_out_pel.full = wr_fifo_mul_9_11_opA.full | wr_fifo_mul_9_18_opA.full | wr_fifo_mul_9_25_opA.full
        | wr_fifo_mul_9_32_opA.full;
        
        // - WRITE 
        assign wr_fifo_mul_9_11_opA.write = wr_delay_3_out_pel.write;
        assign wr_fifo_mul_9_18_opA.write = wr_delay_3_out_pel.write;
        assign wr_fifo_mul_9_25_opA.write = wr_delay_3_out_pel.write;
        assign wr_fifo_mul_9_32_opA.write = wr_delay_3_out_pel.write;
        
        // - DATA
        assign wr_fifo_mul_9_11_opA.din = wr_delay_3_out_pel.din;
        assign wr_fifo_mul_9_18_opA.din = wr_delay_3_out_pel.din;
        assign wr_fifo_mul_9_25_opA.din = wr_delay_3_out_pel.din;
        assign wr_fifo_mul_9_32_opA.din = wr_delay_3_out_pel.din;
    
    //FORK DELAY 4 TO MUL_9_12 & MUL_9_19 & MUL_9_26 & MUL_9_33 & MUL_9_40

        // - INTERFACES   		    		
        write_interface #(8,FLUX) wr_fifo_mul_9_12_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_19_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_26_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_33_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_40_opA(clk);
               
        // - FULL
        assign wr_delay_4_out_pel.full = wr_fifo_mul_9_12_opA.full | wr_fifo_mul_9_19_opA.full | wr_fifo_mul_9_26_opA.full
        | wr_fifo_mul_9_33_opA.full | wr_fifo_mul_9_40_opA.full;
        
        // - WRITE 
        assign wr_fifo_mul_9_12_opA.write = wr_delay_4_out_pel.write;
        assign wr_fifo_mul_9_19_opA.write = wr_delay_4_out_pel.write;
        assign wr_fifo_mul_9_26_opA.write = wr_delay_4_out_pel.write;
        assign wr_fifo_mul_9_33_opA.write = wr_delay_4_out_pel.write;
        assign wr_fifo_mul_9_40_opA.write = wr_delay_4_out_pel.write;
        
        // - DATA
        assign wr_fifo_mul_9_12_opA.din = wr_delay_4_out_pel.din;
        assign wr_fifo_mul_9_19_opA.din = wr_delay_4_out_pel.din;
        assign wr_fifo_mul_9_26_opA.din = wr_delay_4_out_pel.din;
        assign wr_fifo_mul_9_33_opA.din = wr_delay_4_out_pel.din;
        assign wr_fifo_mul_9_40_opA.din = wr_delay_4_out_pel.din;
            
    //FORK DELAY 5 TO MUL_9_13 & MUL_9_20 & MUL_9_27 & MUL_9_34 & MUL_9_41 & MUL_9_48

        // - INTERFACES   		    		
        write_interface #(8,FLUX) wr_fifo_mul_9_13_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_20_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_27_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_34_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_41_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_48_opA(clk); 
               
        // - FULL
        assign wr_delay_5_out_pel.full = wr_fifo_mul_9_13_opA.full | wr_fifo_mul_9_20_opA.full | wr_fifo_mul_9_27_opA.full
        | wr_fifo_mul_9_34_opA.full | wr_fifo_mul_9_41_opA.full | wr_fifo_mul_9_48_opA.full;
        
        // - WRITE 
        assign wr_fifo_mul_9_13_opA.write = wr_delay_5_out_pel.write;
        assign wr_fifo_mul_9_20_opA.write = wr_delay_5_out_pel.write;
        assign wr_fifo_mul_9_27_opA.write = wr_delay_5_out_pel.write;
        assign wr_fifo_mul_9_34_opA.write = wr_delay_5_out_pel.write;
        assign wr_fifo_mul_9_41_opA.write = wr_delay_5_out_pel.write;
        assign wr_fifo_mul_9_48_opA.write = wr_delay_5_out_pel.write;
        
        // - DATA
        assign wr_fifo_mul_9_13_opA.din = wr_delay_5_out_pel.din;
        assign wr_fifo_mul_9_20_opA.din = wr_delay_5_out_pel.din;
        assign wr_fifo_mul_9_27_opA.din = wr_delay_5_out_pel.din;
        assign wr_fifo_mul_9_34_opA.din = wr_delay_5_out_pel.din;
        assign wr_fifo_mul_9_41_opA.din = wr_delay_5_out_pel.din;
        assign wr_fifo_mul_9_48_opA.din = wr_delay_5_out_pel.din;
		
	//FORK DELAY 6 TO MUL_9_14 & MUL_9_21 & MUL_9_28 & MUL_9_35 & MUL_9_42 & MUL_9_49 & MUL_9_56

        // - INTERFACES   		    		
        write_interface #(8,FLUX) wr_fifo_mul_9_14_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_21_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_28_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_35_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_42_opA(clk);
        write_interface #(8,FLUX) wr_fifo_mul_9_49_opA(clk); 
		write_interface #(8,FLUX) wr_fifo_mul_9_56_opA(clk); 
               
        // - FULL
        assign wr_delay_6_out_pel.full = wr_fifo_mul_9_14_opA.full | wr_fifo_mul_9_21_opA.full | wr_fifo_mul_9_28_opA.full
        | wr_fifo_mul_9_35_opA.full | wr_fifo_mul_9_42_opA.full | wr_fifo_mul_9_49_opA.full | wr_fifo_mul_9_56_opA.full;
        
        // - WRITE 
        assign wr_fifo_mul_9_14_opA.write = wr_delay_6_out_pel.write;
        assign wr_fifo_mul_9_21_opA.write = wr_delay_6_out_pel.write;
        assign wr_fifo_mul_9_28_opA.write = wr_delay_6_out_pel.write;
        assign wr_fifo_mul_9_35_opA.write = wr_delay_6_out_pel.write;
        assign wr_fifo_mul_9_42_opA.write = wr_delay_6_out_pel.write;
        assign wr_fifo_mul_9_49_opA.write = wr_delay_6_out_pel.write;
		assign wr_fifo_mul_9_56_opA.write = wr_delay_6_out_pel.write;
        
        // - DATA
        assign wr_fifo_mul_9_14_opA.din = wr_delay_6_out_pel.din;
        assign wr_fifo_mul_9_21_opA.din = wr_delay_6_out_pel.din;
        assign wr_fifo_mul_9_28_opA.din = wr_delay_6_out_pel.din;
        assign wr_fifo_mul_9_35_opA.din = wr_delay_6_out_pel.din;
        assign wr_fifo_mul_9_42_opA.din = wr_delay_6_out_pel.din;
        assign wr_fifo_mul_9_49_opA.din = wr_delay_6_out_pel.din;
		assign wr_fifo_mul_9_56_opA.din = wr_delay_6_out_pel.din;

        
    //FORK coeff h C0 TO MUL_9_0 & MUL_9_8 & MUL_9_16 & MUL_24 & MUL_32 & MUL_40 & MUL_48 & MUL_56
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_9_0_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_8_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_9_16_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_24_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_32_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_40_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_48_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_56_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_h_c0.full = wr_fifo_mul_9_0_opB.full | wr_fifo_mul_9_8_opB.full | wr_fifo_mul_9_16_opB.full 
        | wr_fifo_mul_9_24_opB.full | wr_fifo_mul_9_32_opB.full | wr_fifo_mul_9_40_opB.full | wr_fifo_mul_9_48_opB.full
        | wr_fifo_mul_9_56_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_9_0_opB.write = wr_coeff_luma_h_c0.write;
        assign wr_fifo_mul_9_8_opB.write = wr_coeff_luma_h_c0.write;
        assign wr_fifo_mul_9_16_opB.write = wr_coeff_luma_h_c0.write;
        assign wr_fifo_mul_9_24_opB.write = wr_coeff_luma_h_c0.write;
        assign wr_fifo_mul_9_32_opB.write = wr_coeff_luma_h_c0.write;
        assign wr_fifo_mul_9_40_opB.write = wr_coeff_luma_h_c0.write;
        assign wr_fifo_mul_9_48_opB.write = wr_coeff_luma_h_c0.write;
        assign wr_fifo_mul_9_56_opB.write = wr_coeff_luma_h_c0.write;
        
        // - DATA
        assign wr_fifo_mul_9_0_opB.din = wr_coeff_luma_h_c0.din;
        assign wr_fifo_mul_9_8_opB.din = wr_coeff_luma_h_c0.din;
        assign wr_fifo_mul_9_16_opB.din = wr_coeff_luma_h_c0.din;
        assign wr_fifo_mul_9_24_opB.din = wr_coeff_luma_h_c0.din;
        assign wr_fifo_mul_9_32_opB.din = wr_coeff_luma_h_c0.din;
        assign wr_fifo_mul_9_40_opB.din = wr_coeff_luma_h_c0.din;
        assign wr_fifo_mul_9_48_opB.din = wr_coeff_luma_h_c0.din;
        assign wr_fifo_mul_9_56_opB.din = wr_coeff_luma_h_c0.din;
        
    //FORK coeff h C1 TO MUL_9_1 & MUL_9_9 & MUL_9_17 & MUL_25 & MUL_33 & MUL_41 & MUL_49 & MUL_57
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_9_1_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_9_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_9_17_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_25_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_33_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_41_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_49_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_57_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_h_c1.full = wr_fifo_mul_9_1_opB.full | wr_fifo_mul_9_9_opB.full | wr_fifo_mul_9_17_opB.full 
        | wr_fifo_mul_9_25_opB.full | wr_fifo_mul_9_33_opB.full | wr_fifo_mul_9_41_opB.full | wr_fifo_mul_9_49_opB.full
        | wr_fifo_mul_9_57_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_9_1_opB.write = wr_coeff_luma_h_c1.write;
        assign wr_fifo_mul_9_9_opB.write = wr_coeff_luma_h_c1.write;
        assign wr_fifo_mul_9_17_opB.write = wr_coeff_luma_h_c1.write;
        assign wr_fifo_mul_9_25_opB.write = wr_coeff_luma_h_c1.write;
        assign wr_fifo_mul_9_33_opB.write = wr_coeff_luma_h_c1.write;
        assign wr_fifo_mul_9_41_opB.write = wr_coeff_luma_h_c1.write;
        assign wr_fifo_mul_9_49_opB.write = wr_coeff_luma_h_c1.write;
        assign wr_fifo_mul_9_57_opB.write = wr_coeff_luma_h_c1.write;
        
        // - DATA
        assign wr_fifo_mul_9_1_opB.din = wr_coeff_luma_h_c1.din;
        assign wr_fifo_mul_9_9_opB.din = wr_coeff_luma_h_c1.din;
        assign wr_fifo_mul_9_17_opB.din = wr_coeff_luma_h_c1.din;
        assign wr_fifo_mul_9_25_opB.din = wr_coeff_luma_h_c1.din;
        assign wr_fifo_mul_9_33_opB.din = wr_coeff_luma_h_c1.din;
        assign wr_fifo_mul_9_41_opB.din = wr_coeff_luma_h_c1.din;
        assign wr_fifo_mul_9_49_opB.din = wr_coeff_luma_h_c1.din;
        assign wr_fifo_mul_9_57_opB.din = wr_coeff_luma_h_c1.din;            
    
    //FORK coeff h C2 TO MUL_9_2 & MUL_9_10 & MUL_9_18 & MUL_26 & MUL_34 & MUL_42 & MUL_50 & MUL_58
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_9_2_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_10_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_9_18_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_26_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_34_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_42_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_50_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_58_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_h_c2.full = wr_fifo_mul_9_2_opB.full | wr_fifo_mul_9_10_opB.full | wr_fifo_mul_9_18_opB.full 
        | wr_fifo_mul_9_26_opB.full | wr_fifo_mul_9_34_opB.full | wr_fifo_mul_9_42_opB.full | wr_fifo_mul_9_50_opB.full
        | wr_fifo_mul_9_58_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_9_2_opB.write = wr_coeff_luma_h_c2.write;
        assign wr_fifo_mul_9_10_opB.write = wr_coeff_luma_h_c2.write;
        assign wr_fifo_mul_9_18_opB.write = wr_coeff_luma_h_c2.write;
        assign wr_fifo_mul_9_26_opB.write = wr_coeff_luma_h_c2.write;
        assign wr_fifo_mul_9_34_opB.write = wr_coeff_luma_h_c2.write;
        assign wr_fifo_mul_9_42_opB.write = wr_coeff_luma_h_c2.write;
        assign wr_fifo_mul_9_50_opB.write = wr_coeff_luma_h_c2.write;
        assign wr_fifo_mul_9_58_opB.write = wr_coeff_luma_h_c2.write;
        
        // - DATA
        assign wr_fifo_mul_9_2_opB.din = wr_coeff_luma_h_c2.din;
        assign wr_fifo_mul_9_10_opB.din = wr_coeff_luma_h_c2.din;
        assign wr_fifo_mul_9_18_opB.din = wr_coeff_luma_h_c2.din;
        assign wr_fifo_mul_9_26_opB.din = wr_coeff_luma_h_c2.din;
        assign wr_fifo_mul_9_34_opB.din = wr_coeff_luma_h_c2.din;
        assign wr_fifo_mul_9_42_opB.din = wr_coeff_luma_h_c2.din;
        assign wr_fifo_mul_9_50_opB.din = wr_coeff_luma_h_c2.din;
        assign wr_fifo_mul_9_58_opB.din = wr_coeff_luma_h_c2.din;
        
    //FORK coeff h C3 TO MUL_9_3 & MUL_9_11 & MUL_9_19 & MUL_27 & MUL_35 & MUL_43 & MUL_51 & MUL_59
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_9_3_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_11_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_9_19_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_27_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_35_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_43_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_51_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_59_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_h_c3.full = wr_fifo_mul_9_3_opB.full | wr_fifo_mul_9_11_opB.full | wr_fifo_mul_9_19_opB.full 
        | wr_fifo_mul_9_27_opB.full | wr_fifo_mul_9_35_opB.full | wr_fifo_mul_9_43_opB.full | wr_fifo_mul_9_51_opB.full
        | wr_fifo_mul_9_59_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_9_3_opB.write = wr_coeff_luma_h_c3.write;
        assign wr_fifo_mul_9_11_opB.write = wr_coeff_luma_h_c3.write;
        assign wr_fifo_mul_9_19_opB.write = wr_coeff_luma_h_c3.write;
        assign wr_fifo_mul_9_27_opB.write = wr_coeff_luma_h_c3.write;
        assign wr_fifo_mul_9_35_opB.write = wr_coeff_luma_h_c3.write;
        assign wr_fifo_mul_9_43_opB.write = wr_coeff_luma_h_c3.write;
        assign wr_fifo_mul_9_51_opB.write = wr_coeff_luma_h_c3.write;
        assign wr_fifo_mul_9_59_opB.write = wr_coeff_luma_h_c3.write;
        
        // - DATA
        assign wr_fifo_mul_9_3_opB.din = wr_coeff_luma_h_c3.din;
        assign wr_fifo_mul_9_11_opB.din = wr_coeff_luma_h_c3.din;
        assign wr_fifo_mul_9_19_opB.din = wr_coeff_luma_h_c3.din;
        assign wr_fifo_mul_9_27_opB.din = wr_coeff_luma_h_c3.din;
        assign wr_fifo_mul_9_35_opB.din = wr_coeff_luma_h_c3.din;
        assign wr_fifo_mul_9_43_opB.din = wr_coeff_luma_h_c3.din;
        assign wr_fifo_mul_9_51_opB.din = wr_coeff_luma_h_c3.din;
        assign wr_fifo_mul_9_59_opB.din = wr_coeff_luma_h_c3.din;        

    //FORK coeff h C4 TO MUL_9_4 & MUL_9_12 & MUL_9_20 & MUL_28 & MUL_36 & MUL_44 & MUL_52 & MUL_60
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_9_4_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_12_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_9_20_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_28_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_36_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_44_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_52_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_60_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_h_c4.full = wr_fifo_mul_9_4_opB.full | wr_fifo_mul_9_12_opB.full | wr_fifo_mul_9_20_opB.full 
        | wr_fifo_mul_9_28_opB.full | wr_fifo_mul_9_36_opB.full | wr_fifo_mul_9_44_opB.full | wr_fifo_mul_9_52_opB.full
        | wr_fifo_mul_9_60_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_9_4_opB.write = wr_coeff_luma_h_c4.write;
        assign wr_fifo_mul_9_12_opB.write = wr_coeff_luma_h_c4.write;
        assign wr_fifo_mul_9_20_opB.write = wr_coeff_luma_h_c4.write;
        assign wr_fifo_mul_9_28_opB.write = wr_coeff_luma_h_c4.write;
        assign wr_fifo_mul_9_36_opB.write = wr_coeff_luma_h_c4.write;
        assign wr_fifo_mul_9_44_opB.write = wr_coeff_luma_h_c4.write;
        assign wr_fifo_mul_9_52_opB.write = wr_coeff_luma_h_c4.write;
        assign wr_fifo_mul_9_60_opB.write = wr_coeff_luma_h_c4.write;
        
        // - DATA
        assign wr_fifo_mul_9_4_opB.din = wr_coeff_luma_h_c4.din;
        assign wr_fifo_mul_9_12_opB.din = wr_coeff_luma_h_c4.din;
        assign wr_fifo_mul_9_20_opB.din = wr_coeff_luma_h_c4.din;
        assign wr_fifo_mul_9_28_opB.din = wr_coeff_luma_h_c4.din;
        assign wr_fifo_mul_9_36_opB.din = wr_coeff_luma_h_c4.din;
        assign wr_fifo_mul_9_44_opB.din = wr_coeff_luma_h_c4.din;
        assign wr_fifo_mul_9_52_opB.din = wr_coeff_luma_h_c4.din;
        assign wr_fifo_mul_9_60_opB.din = wr_coeff_luma_h_c4.din;

    //FORK coeff h C5 TO MUL_9_5 & MUL_9_13 & MUL_9_21 & MUL_29 & MUL_37 & MUL_45 & MUL_53 & MUL_61
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_9_5_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_13_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_9_21_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_29_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_37_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_45_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_53_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_61_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_h_c5.full = wr_fifo_mul_9_5_opB.full | wr_fifo_mul_9_13_opB.full | wr_fifo_mul_9_21_opB.full 
        | wr_fifo_mul_9_29_opB.full | wr_fifo_mul_9_37_opB.full | wr_fifo_mul_9_45_opB.full | wr_fifo_mul_9_53_opB.full
        | wr_fifo_mul_9_61_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_9_5_opB.write = wr_coeff_luma_h_c5.write;
        assign wr_fifo_mul_9_13_opB.write = wr_coeff_luma_h_c5.write;
        assign wr_fifo_mul_9_21_opB.write = wr_coeff_luma_h_c5.write;
        assign wr_fifo_mul_9_29_opB.write = wr_coeff_luma_h_c5.write;
        assign wr_fifo_mul_9_37_opB.write = wr_coeff_luma_h_c5.write;
        assign wr_fifo_mul_9_45_opB.write = wr_coeff_luma_h_c5.write;
        assign wr_fifo_mul_9_53_opB.write = wr_coeff_luma_h_c5.write;
        assign wr_fifo_mul_9_61_opB.write = wr_coeff_luma_h_c5.write;
        
        // - DATA
        assign wr_fifo_mul_9_5_opB.din = wr_coeff_luma_h_c5.din;
        assign wr_fifo_mul_9_13_opB.din = wr_coeff_luma_h_c5.din;
        assign wr_fifo_mul_9_21_opB.din = wr_coeff_luma_h_c5.din;
        assign wr_fifo_mul_9_29_opB.din = wr_coeff_luma_h_c5.din;
        assign wr_fifo_mul_9_37_opB.din = wr_coeff_luma_h_c5.din;
        assign wr_fifo_mul_9_45_opB.din = wr_coeff_luma_h_c5.din;
        assign wr_fifo_mul_9_53_opB.din = wr_coeff_luma_h_c5.din;
        assign wr_fifo_mul_9_61_opB.din = wr_coeff_luma_h_c5.din;
        
    //FORK coeff h C6 TO MUL_9_6 & MUL_9_14 & MUL_9_22 & MUL_30 & MUL_38 & MUL_46 & MUL_54 & MUL_62
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_9_6_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_14_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_9_22_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_30_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_38_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_46_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_54_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_62_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_h_c6.full = wr_fifo_mul_9_6_opB.full | wr_fifo_mul_9_14_opB.full | wr_fifo_mul_9_22_opB.full 
        | wr_fifo_mul_9_30_opB.full | wr_fifo_mul_9_38_opB.full | wr_fifo_mul_9_46_opB.full | wr_fifo_mul_9_54_opB.full
        | wr_fifo_mul_9_62_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_9_6_opB.write = wr_coeff_luma_h_c6.write;
        assign wr_fifo_mul_9_14_opB.write = wr_coeff_luma_h_c6.write;
        assign wr_fifo_mul_9_22_opB.write = wr_coeff_luma_h_c6.write;
        assign wr_fifo_mul_9_30_opB.write = wr_coeff_luma_h_c6.write;
        assign wr_fifo_mul_9_38_opB.write = wr_coeff_luma_h_c6.write;
        assign wr_fifo_mul_9_46_opB.write = wr_coeff_luma_h_c6.write;
        assign wr_fifo_mul_9_54_opB.write = wr_coeff_luma_h_c6.write;
        assign wr_fifo_mul_9_62_opB.write = wr_coeff_luma_h_c6.write;
        
        // - DATA
        assign wr_fifo_mul_9_6_opB.din = wr_coeff_luma_h_c6.din;
        assign wr_fifo_mul_9_14_opB.din = wr_coeff_luma_h_c6.din;
        assign wr_fifo_mul_9_22_opB.din = wr_coeff_luma_h_c6.din;
        assign wr_fifo_mul_9_30_opB.din = wr_coeff_luma_h_c6.din;
        assign wr_fifo_mul_9_38_opB.din = wr_coeff_luma_h_c6.din;
        assign wr_fifo_mul_9_46_opB.din = wr_coeff_luma_h_c6.din;
        assign wr_fifo_mul_9_54_opB.din = wr_coeff_luma_h_c6.din;
        assign wr_fifo_mul_9_62_opB.din = wr_coeff_luma_h_c6.din;        

    //FORK coeff h C7 TO MUL_9_7 & MUL_9_15 & MUL_9_23 & MUL_31 & MUL_39 & MUL_47 & MUL_55 & MUL_63
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_9_7_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_15_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_9_23_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_31_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_39_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_47_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_55_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_9_63_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_h_c7.full = wr_fifo_mul_9_7_opB.full | wr_fifo_mul_9_15_opB.full | wr_fifo_mul_9_23_opB.full 
        | wr_fifo_mul_9_31_opB.full | wr_fifo_mul_9_39_opB.full | wr_fifo_mul_9_47_opB.full | wr_fifo_mul_9_55_opB.full
        | wr_fifo_mul_9_63_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_9_7_opB.write = wr_coeff_luma_h_c7.write;
        assign wr_fifo_mul_9_15_opB.write = wr_coeff_luma_h_c7.write;
        assign wr_fifo_mul_9_23_opB.write = wr_coeff_luma_h_c7.write;
        assign wr_fifo_mul_9_31_opB.write = wr_coeff_luma_h_c7.write;
        assign wr_fifo_mul_9_39_opB.write = wr_coeff_luma_h_c7.write;
        assign wr_fifo_mul_9_47_opB.write = wr_coeff_luma_h_c7.write;
        assign wr_fifo_mul_9_55_opB.write = wr_coeff_luma_h_c7.write;
        assign wr_fifo_mul_9_63_opB.write = wr_coeff_luma_h_c7.write;
        
        // - DATA
        assign wr_fifo_mul_9_7_opB.din = wr_coeff_luma_h_c7.din;
        assign wr_fifo_mul_9_15_opB.din = wr_coeff_luma_h_c7.din;
        assign wr_fifo_mul_9_23_opB.din = wr_coeff_luma_h_c7.din;
        assign wr_fifo_mul_9_31_opB.din = wr_coeff_luma_h_c7.din;
        assign wr_fifo_mul_9_39_opB.din = wr_coeff_luma_h_c7.din;
        assign wr_fifo_mul_9_47_opB.din = wr_coeff_luma_h_c7.din;
        assign wr_fifo_mul_9_55_opB.din = wr_coeff_luma_h_c7.din;
        assign wr_fifo_mul_9_63_opB.din = wr_coeff_luma_h_c7.din;
 
        
    //FORKS SECONDA PARTE
    
    //FORK REMOVE_h to mul_18_0 & mul_18_8 & mul_18_16 & mul_18_24 & mul_18_32 & mul_18_40 & mul_18_48 & mul_18_56
    
        // - INTERFACES 
        write_interface #(18,FLUX) wr_fifo_line_buffer_0_0_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_0_1_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_0_2_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_0_3_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_0_4_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_0_5_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_0_6_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_0_7_in_pel(clk);
        
        write_interface #(18,FLUX) wr_fifo_mul_18_0_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_8_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_16_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_24_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_32_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_40_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_48_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_56_opA(clk);               
     
        // - FULL
        assign wr_remove_h_0_out_pel.full = wr_fifo_line_buffer_0_0_in_pel.full | wr_fifo_mul_18_0_opA.full;
        assign wr_remove_h_1_out_pel.full = wr_fifo_line_buffer_0_1_in_pel.full | wr_fifo_mul_18_8_opA.full;
        assign wr_remove_h_2_out_pel.full = wr_fifo_line_buffer_0_2_in_pel.full | wr_fifo_mul_18_16_opA.full;
        assign wr_remove_h_3_out_pel.full = wr_fifo_line_buffer_0_3_in_pel.full | wr_fifo_mul_18_24_opA.full;
        assign wr_remove_h_4_out_pel.full = wr_fifo_line_buffer_0_4_in_pel.full | wr_fifo_mul_18_32_opA.full;
        assign wr_remove_h_5_out_pel.full = wr_fifo_line_buffer_0_5_in_pel.full | wr_fifo_mul_18_40_opA.full;
        assign wr_remove_h_6_out_pel.full = wr_fifo_line_buffer_0_6_in_pel.full | wr_fifo_mul_18_48_opA.full;
        assign wr_remove_h_7_out_pel.full = wr_fifo_line_buffer_0_7_in_pel.full | wr_fifo_mul_18_56_opA.full;
     
        // - WRITE
        assign wr_fifo_line_buffer_0_0_in_pel.write = wr_remove_h_0_out_pel.write;
        assign wr_fifo_mul_18_0_opA.write = wr_remove_h_0_out_pel.write;
        assign wr_fifo_line_buffer_0_1_in_pel.write = wr_remove_h_1_out_pel.write;
        assign wr_fifo_mul_18_8_opA.write = wr_remove_h_1_out_pel.write;
        assign wr_fifo_line_buffer_0_2_in_pel.write = wr_remove_h_2_out_pel.write;
        assign wr_fifo_mul_18_16_opA.write = wr_remove_h_2_out_pel.write;     
        assign wr_fifo_line_buffer_0_3_in_pel.write = wr_remove_h_3_out_pel.write;
        assign wr_fifo_mul_18_24_opA.write = wr_remove_h_3_out_pel.write;
        assign wr_fifo_line_buffer_0_4_in_pel.write = wr_remove_h_4_out_pel.write;
        assign wr_fifo_mul_18_32_opA.write = wr_remove_h_4_out_pel.write;     
        assign wr_fifo_line_buffer_0_5_in_pel.write = wr_remove_h_5_out_pel.write;
        assign wr_fifo_mul_18_40_opA.write = wr_remove_h_5_out_pel.write;
        assign wr_fifo_line_buffer_0_6_in_pel.write = wr_remove_h_6_out_pel.write;
        assign wr_fifo_mul_18_48_opA.write = wr_remove_h_6_out_pel.write;     
        assign wr_fifo_line_buffer_0_7_in_pel.write = wr_remove_h_7_out_pel.write;
        assign wr_fifo_mul_18_56_opA.write = wr_remove_h_7_out_pel.write;
                        
        // - DATA
        assign wr_fifo_line_buffer_0_0_in_pel.din = wr_remove_h_0_out_pel.din;
        assign wr_fifo_mul_18_0_opA.din = wr_remove_h_0_out_pel.din;
        assign wr_fifo_line_buffer_0_1_in_pel.din = wr_remove_h_1_out_pel.din;
        assign wr_fifo_mul_18_8_opA.din = wr_remove_h_1_out_pel.din;
        assign wr_fifo_line_buffer_0_2_in_pel.din = wr_remove_h_2_out_pel.din;
        assign wr_fifo_mul_18_16_opA.din = wr_remove_h_2_out_pel.din;     
        assign wr_fifo_line_buffer_0_3_in_pel.din = wr_remove_h_3_out_pel.din;
        assign wr_fifo_mul_18_24_opA.din = wr_remove_h_3_out_pel.din;
        assign wr_fifo_line_buffer_0_4_in_pel.din = wr_remove_h_4_out_pel.din;
        assign wr_fifo_mul_18_32_opA.din = wr_remove_h_4_out_pel.din;     
        assign wr_fifo_line_buffer_0_5_in_pel.din = wr_remove_h_5_out_pel.din;
        assign wr_fifo_mul_18_40_opA.din = wr_remove_h_5_out_pel.din;
        assign wr_fifo_line_buffer_0_6_in_pel.din = wr_remove_h_6_out_pel.din;
        assign wr_fifo_mul_18_48_opA.din = wr_remove_h_6_out_pel.din;     
        assign wr_fifo_line_buffer_0_7_in_pel.din = wr_remove_h_7_out_pel.din;
        assign wr_fifo_mul_18_56_opA.din = wr_remove_h_7_out_pel.din;    
    
    //FORK line_buffer_0 to mul_18_1 & mul_18_9 & mul_18_17 & mul_18_25 & mul_18_33 & mul_18_41 & mul_18_49 & mul_18_57
    
        // - INTERFACES 
        write_interface #(18,FLUX) wr_fifo_line_buffer_1_0_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_1_1_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_1_2_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_1_3_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_1_4_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_1_5_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_1_6_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_1_7_in_pel(clk);
        
        write_interface #(18,FLUX) wr_fifo_mul_18_1_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_9_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_17_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_25_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_33_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_41_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_49_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_57_opA(clk);               
     
        // - FULL
        assign wr_line_buffer_0_0_out_pel.full = wr_fifo_line_buffer_1_0_in_pel.full | wr_fifo_mul_18_1_opA.full;
        assign wr_line_buffer_0_1_out_pel.full = wr_fifo_line_buffer_1_1_in_pel.full | wr_fifo_mul_18_9_opA.full;
        assign wr_line_buffer_0_2_out_pel.full = wr_fifo_line_buffer_1_2_in_pel.full | wr_fifo_mul_18_17_opA.full;
        assign wr_line_buffer_0_3_out_pel.full = wr_fifo_line_buffer_1_3_in_pel.full | wr_fifo_mul_18_25_opA.full;
        assign wr_line_buffer_0_4_out_pel.full = wr_fifo_line_buffer_1_4_in_pel.full | wr_fifo_mul_18_33_opA.full;
        assign wr_line_buffer_0_5_out_pel.full = wr_fifo_line_buffer_1_5_in_pel.full | wr_fifo_mul_18_41_opA.full;
        assign wr_line_buffer_0_6_out_pel.full = wr_fifo_line_buffer_1_6_in_pel.full | wr_fifo_mul_18_49_opA.full;
        assign wr_line_buffer_0_7_out_pel.full = wr_fifo_line_buffer_1_7_in_pel.full | wr_fifo_mul_18_57_opA.full;
     
        // - WRITE
        assign wr_fifo_line_buffer_1_0_in_pel.write = wr_line_buffer_0_0_out_pel.write;
        assign wr_fifo_mul_18_1_opA.write = wr_line_buffer_0_0_out_pel.write;
        assign wr_fifo_line_buffer_1_1_in_pel.write = wr_line_buffer_0_1_out_pel.write;
        assign wr_fifo_mul_18_9_opA.write = wr_line_buffer_0_1_out_pel.write;
        assign wr_fifo_line_buffer_1_2_in_pel.write = wr_line_buffer_0_2_out_pel.write;
        assign wr_fifo_mul_18_17_opA.write = wr_line_buffer_0_2_out_pel.write;     
        assign wr_fifo_line_buffer_1_3_in_pel.write = wr_line_buffer_0_3_out_pel.write;
        assign wr_fifo_mul_18_25_opA.write = wr_line_buffer_0_3_out_pel.write;
        assign wr_fifo_line_buffer_1_4_in_pel.write = wr_line_buffer_0_4_out_pel.write;
        assign wr_fifo_mul_18_33_opA.write = wr_line_buffer_0_4_out_pel.write;     
        assign wr_fifo_line_buffer_1_5_in_pel.write = wr_line_buffer_0_5_out_pel.write;
        assign wr_fifo_mul_18_41_opA.write = wr_line_buffer_0_5_out_pel.write;
        assign wr_fifo_line_buffer_1_6_in_pel.write = wr_line_buffer_0_6_out_pel.write;
        assign wr_fifo_mul_18_49_opA.write = wr_line_buffer_0_6_out_pel.write;     
        assign wr_fifo_line_buffer_1_7_in_pel.write = wr_line_buffer_0_7_out_pel.write;
        assign wr_fifo_mul_18_57_opA.write = wr_line_buffer_0_7_out_pel.write;
                        
        // - DATA
        assign wr_fifo_line_buffer_1_0_in_pel.din = wr_line_buffer_0_0_out_pel.din;
        assign wr_fifo_mul_18_1_opA.din = wr_line_buffer_0_0_out_pel.din;
        assign wr_fifo_line_buffer_1_1_in_pel.din = wr_line_buffer_0_1_out_pel.din;
        assign wr_fifo_mul_18_9_opA.din = wr_line_buffer_0_1_out_pel.din;
        assign wr_fifo_line_buffer_1_2_in_pel.din = wr_line_buffer_0_2_out_pel.din;
        assign wr_fifo_mul_18_17_opA.din = wr_line_buffer_0_2_out_pel.din;     
        assign wr_fifo_line_buffer_1_3_in_pel.din = wr_line_buffer_0_3_out_pel.din;
        assign wr_fifo_mul_18_25_opA.din = wr_line_buffer_0_3_out_pel.din;
        assign wr_fifo_line_buffer_1_4_in_pel.din = wr_line_buffer_0_4_out_pel.din;
        assign wr_fifo_mul_18_33_opA.din = wr_line_buffer_0_4_out_pel.din;     
        assign wr_fifo_line_buffer_1_5_in_pel.din = wr_line_buffer_0_5_out_pel.din;
        assign wr_fifo_mul_18_41_opA.din = wr_line_buffer_0_5_out_pel.din;
        assign wr_fifo_line_buffer_1_6_in_pel.din = wr_line_buffer_0_6_out_pel.din;
        assign wr_fifo_mul_18_49_opA.din = wr_line_buffer_0_6_out_pel.din;     
        assign wr_fifo_line_buffer_1_7_in_pel.din = wr_line_buffer_0_7_out_pel.din;
        assign wr_fifo_mul_18_57_opA.din = wr_line_buffer_0_7_out_pel.din;
        
    //FORK line_buffer_1 to mul_18_2 & mul_18_10 & mul_18_18 & mul_18_26 & mul_18_34 & mul_18_42 & mul_18_50 & mul_18_58
    
        // - INTERFACES 
        write_interface #(18,FLUX) wr_fifo_line_buffer_2_0_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_2_1_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_2_2_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_2_3_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_2_4_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_2_5_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_2_6_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_2_7_in_pel(clk);    

        write_interface #(18,FLUX) wr_fifo_mul_18_2_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_10_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_18_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_26_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_34_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_42_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_50_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_58_opA(clk);               
     
        // - FULL
        assign wr_line_buffer_1_0_out_pel.full = wr_fifo_line_buffer_2_0_in_pel.full | wr_fifo_mul_18_2_opA.full;
        assign wr_line_buffer_1_1_out_pel.full = wr_fifo_line_buffer_2_1_in_pel.full | wr_fifo_mul_18_10_opA.full;
        assign wr_line_buffer_1_2_out_pel.full = wr_fifo_line_buffer_2_2_in_pel.full | wr_fifo_mul_18_18_opA.full;
        assign wr_line_buffer_1_3_out_pel.full = wr_fifo_line_buffer_2_3_in_pel.full | wr_fifo_mul_18_26_opA.full;
        assign wr_line_buffer_1_4_out_pel.full = wr_fifo_line_buffer_2_4_in_pel.full | wr_fifo_mul_18_34_opA.full;
        assign wr_line_buffer_1_5_out_pel.full = wr_fifo_line_buffer_2_5_in_pel.full | wr_fifo_mul_18_42_opA.full;
        assign wr_line_buffer_1_6_out_pel.full = wr_fifo_line_buffer_2_6_in_pel.full | wr_fifo_mul_18_50_opA.full;
        assign wr_line_buffer_1_7_out_pel.full = wr_fifo_line_buffer_2_7_in_pel.full | wr_fifo_mul_18_58_opA.full;
     
        // - WRITE
        assign wr_fifo_line_buffer_2_0_in_pel.write = wr_line_buffer_1_0_out_pel.write;
        assign wr_fifo_mul_18_2_opA.write = wr_line_buffer_1_0_out_pel.write;
        assign wr_fifo_line_buffer_2_1_in_pel.write = wr_line_buffer_1_1_out_pel.write;
        assign wr_fifo_mul_18_10_opA.write = wr_line_buffer_1_1_out_pel.write;
        assign wr_fifo_line_buffer_2_2_in_pel.write = wr_line_buffer_1_2_out_pel.write;
        assign wr_fifo_mul_18_18_opA.write = wr_line_buffer_1_2_out_pel.write;     
        assign wr_fifo_line_buffer_2_3_in_pel.write = wr_line_buffer_1_3_out_pel.write;
        assign wr_fifo_mul_18_26_opA.write = wr_line_buffer_1_3_out_pel.write;
        assign wr_fifo_line_buffer_2_4_in_pel.write = wr_line_buffer_1_4_out_pel.write;
        assign wr_fifo_mul_18_34_opA.write = wr_line_buffer_1_4_out_pel.write;     
        assign wr_fifo_line_buffer_2_5_in_pel.write = wr_line_buffer_1_5_out_pel.write;
        assign wr_fifo_mul_18_42_opA.write = wr_line_buffer_1_5_out_pel.write;
        assign wr_fifo_line_buffer_2_6_in_pel.write = wr_line_buffer_1_6_out_pel.write;
        assign wr_fifo_mul_18_50_opA.write = wr_line_buffer_1_6_out_pel.write;     
        assign wr_fifo_line_buffer_2_7_in_pel.write = wr_line_buffer_1_7_out_pel.write;
        assign wr_fifo_mul_18_58_opA.write = wr_line_buffer_1_7_out_pel.write;
                        
        // - DATA
        assign wr_fifo_line_buffer_2_0_in_pel.din = wr_line_buffer_1_0_out_pel.din;
        assign wr_fifo_mul_18_2_opA.din = wr_line_buffer_1_0_out_pel.din;
        assign wr_fifo_line_buffer_2_1_in_pel.din = wr_line_buffer_1_1_out_pel.din;
        assign wr_fifo_mul_18_10_opA.din = wr_line_buffer_1_1_out_pel.din;
        assign wr_fifo_line_buffer_2_2_in_pel.din = wr_line_buffer_1_2_out_pel.din;
        assign wr_fifo_mul_18_18_opA.din = wr_line_buffer_1_2_out_pel.din;     
        assign wr_fifo_line_buffer_2_3_in_pel.din = wr_line_buffer_1_3_out_pel.din;
        assign wr_fifo_mul_18_26_opA.din = wr_line_buffer_1_3_out_pel.din;
        assign wr_fifo_line_buffer_2_4_in_pel.din = wr_line_buffer_1_4_out_pel.din;
        assign wr_fifo_mul_18_34_opA.din = wr_line_buffer_1_4_out_pel.din;     
        assign wr_fifo_line_buffer_2_5_in_pel.din = wr_line_buffer_1_5_out_pel.din;
        assign wr_fifo_mul_18_42_opA.din = wr_line_buffer_1_5_out_pel.din;
        assign wr_fifo_line_buffer_2_6_in_pel.din = wr_line_buffer_1_6_out_pel.din;
        assign wr_fifo_mul_18_50_opA.din = wr_line_buffer_1_6_out_pel.din;     
        assign wr_fifo_line_buffer_2_7_in_pel.din = wr_line_buffer_1_7_out_pel.din;
        assign wr_fifo_mul_18_58_opA.din = wr_line_buffer_1_7_out_pel.din;
    
    //FORK line_buffer_2 to mul_18_3 & mul_18_11 & mul_18_19 & mul_18_27 & mul_18_35 & mul_18_43 & mul_18_51 & mul_18_59

        // - INTERFACES 
        write_interface #(18,FLUX) wr_fifo_line_buffer_3_0_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_3_1_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_3_2_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_3_3_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_3_4_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_3_5_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_3_6_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_3_7_in_pel(clk);
        
        write_interface #(18,FLUX) wr_fifo_mul_18_3_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_11_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_19_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_27_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_35_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_43_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_51_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_59_opA(clk);               
     
        // - FULL
        assign wr_line_buffer_2_0_out_pel.full = wr_fifo_line_buffer_3_0_in_pel.full | wr_fifo_mul_18_3_opA.full;
        assign wr_line_buffer_2_1_out_pel.full = wr_fifo_line_buffer_3_1_in_pel.full | wr_fifo_mul_18_11_opA.full;
        assign wr_line_buffer_2_2_out_pel.full = wr_fifo_line_buffer_3_2_in_pel.full | wr_fifo_mul_18_19_opA.full;
        assign wr_line_buffer_2_3_out_pel.full = wr_fifo_line_buffer_3_3_in_pel.full | wr_fifo_mul_18_27_opA.full;
        assign wr_line_buffer_2_4_out_pel.full = wr_fifo_line_buffer_3_4_in_pel.full | wr_fifo_mul_18_35_opA.full;
        assign wr_line_buffer_2_5_out_pel.full = wr_fifo_line_buffer_3_5_in_pel.full | wr_fifo_mul_18_43_opA.full;
        assign wr_line_buffer_2_6_out_pel.full = wr_fifo_line_buffer_3_6_in_pel.full | wr_fifo_mul_18_51_opA.full;
        assign wr_line_buffer_2_7_out_pel.full = wr_fifo_line_buffer_3_7_in_pel.full | wr_fifo_mul_18_59_opA.full;
     
        // - WRITE
        assign wr_fifo_line_buffer_3_0_in_pel.write = wr_line_buffer_2_0_out_pel.write;
        assign wr_fifo_mul_18_3_opA.write = wr_line_buffer_2_0_out_pel.write;
        assign wr_fifo_line_buffer_3_1_in_pel.write = wr_line_buffer_2_1_out_pel.write;
        assign wr_fifo_mul_18_11_opA.write = wr_line_buffer_2_1_out_pel.write;
        assign wr_fifo_line_buffer_3_2_in_pel.write = wr_line_buffer_2_2_out_pel.write;
        assign wr_fifo_mul_18_19_opA.write = wr_line_buffer_2_2_out_pel.write;     
        assign wr_fifo_line_buffer_3_3_in_pel.write = wr_line_buffer_2_3_out_pel.write;
        assign wr_fifo_mul_18_27_opA.write = wr_line_buffer_2_3_out_pel.write;
        assign wr_fifo_line_buffer_3_4_in_pel.write = wr_line_buffer_2_4_out_pel.write;
        assign wr_fifo_mul_18_35_opA.write = wr_line_buffer_2_4_out_pel.write;     
        assign wr_fifo_line_buffer_3_5_in_pel.write = wr_line_buffer_2_5_out_pel.write;
        assign wr_fifo_mul_18_43_opA.write = wr_line_buffer_2_5_out_pel.write;
        assign wr_fifo_line_buffer_3_6_in_pel.write = wr_line_buffer_2_6_out_pel.write;
        assign wr_fifo_mul_18_51_opA.write = wr_line_buffer_2_6_out_pel.write;     
        assign wr_fifo_line_buffer_3_7_in_pel.write = wr_line_buffer_2_7_out_pel.write;
        assign wr_fifo_mul_18_59_opA.write = wr_line_buffer_2_7_out_pel.write;
                        
        // - DATA
        assign wr_fifo_line_buffer_3_0_in_pel.din = wr_line_buffer_2_0_out_pel.din;
        assign wr_fifo_mul_18_3_opA.din = wr_line_buffer_2_0_out_pel.din;
        assign wr_fifo_line_buffer_3_1_in_pel.din = wr_line_buffer_2_1_out_pel.din;
        assign wr_fifo_mul_18_11_opA.din = wr_line_buffer_2_1_out_pel.din;
        assign wr_fifo_line_buffer_3_2_in_pel.din = wr_line_buffer_2_2_out_pel.din;
        assign wr_fifo_mul_18_19_opA.din = wr_line_buffer_2_2_out_pel.din;     
        assign wr_fifo_line_buffer_3_3_in_pel.din = wr_line_buffer_2_3_out_pel.din;
        assign wr_fifo_mul_18_27_opA.din = wr_line_buffer_2_3_out_pel.din;
        assign wr_fifo_line_buffer_3_4_in_pel.din = wr_line_buffer_2_4_out_pel.din;
        assign wr_fifo_mul_18_35_opA.din = wr_line_buffer_2_4_out_pel.din;     
        assign wr_fifo_line_buffer_3_5_in_pel.din = wr_line_buffer_2_5_out_pel.din;
        assign wr_fifo_mul_18_43_opA.din = wr_line_buffer_2_5_out_pel.din;
        assign wr_fifo_line_buffer_3_6_in_pel.din = wr_line_buffer_2_6_out_pel.din;
        assign wr_fifo_mul_18_51_opA.din = wr_line_buffer_2_6_out_pel.din;     
        assign wr_fifo_line_buffer_3_7_in_pel.din = wr_line_buffer_2_7_out_pel.din;
        assign wr_fifo_mul_18_59_opA.din = wr_line_buffer_2_7_out_pel.din;
    
    //FORK line_buffer_3 to mul_18_4 & mul_18_12 & mul_18_20 & mul_18_28 & mul_18_36 & mul_18_44 & mul_18_52 & mul_18_60

        // - INTERFACES 
        write_interface #(18,FLUX) wr_fifo_line_buffer_4_0_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_4_1_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_4_2_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_4_3_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_4_4_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_4_5_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_4_6_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_4_7_in_pel(clk);
        
        write_interface #(18,FLUX) wr_fifo_mul_18_4_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_12_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_20_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_28_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_36_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_44_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_52_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_60_opA(clk);               
     
        // - FULL
        assign wr_line_buffer_3_0_out_pel.full = wr_fifo_line_buffer_4_0_in_pel.full | wr_fifo_mul_18_4_opA.full;
        assign wr_line_buffer_3_1_out_pel.full = wr_fifo_line_buffer_4_1_in_pel.full | wr_fifo_mul_18_12_opA.full;
        assign wr_line_buffer_3_2_out_pel.full = wr_fifo_line_buffer_4_2_in_pel.full | wr_fifo_mul_18_20_opA.full;
        assign wr_line_buffer_3_3_out_pel.full = wr_fifo_line_buffer_4_3_in_pel.full | wr_fifo_mul_18_28_opA.full;
        assign wr_line_buffer_3_4_out_pel.full = wr_fifo_line_buffer_4_4_in_pel.full | wr_fifo_mul_18_36_opA.full;
        assign wr_line_buffer_3_5_out_pel.full = wr_fifo_line_buffer_4_5_in_pel.full | wr_fifo_mul_18_44_opA.full;
        assign wr_line_buffer_3_6_out_pel.full = wr_fifo_line_buffer_4_6_in_pel.full | wr_fifo_mul_18_52_opA.full;
        assign wr_line_buffer_3_7_out_pel.full = wr_fifo_line_buffer_4_7_in_pel.full | wr_fifo_mul_18_60_opA.full;
     
        // - WRITE
        assign wr_fifo_line_buffer_4_0_in_pel.write = wr_line_buffer_3_0_out_pel.write;
        assign wr_fifo_mul_18_4_opA.write = wr_line_buffer_3_0_out_pel.write;
        assign wr_fifo_line_buffer_4_1_in_pel.write = wr_line_buffer_3_1_out_pel.write;
        assign wr_fifo_mul_18_12_opA.write = wr_line_buffer_3_1_out_pel.write;
        assign wr_fifo_line_buffer_4_2_in_pel.write = wr_line_buffer_3_2_out_pel.write;
        assign wr_fifo_mul_18_20_opA.write = wr_line_buffer_3_2_out_pel.write;     
        assign wr_fifo_line_buffer_4_3_in_pel.write = wr_line_buffer_3_3_out_pel.write;
        assign wr_fifo_mul_18_28_opA.write = wr_line_buffer_3_3_out_pel.write;
        assign wr_fifo_line_buffer_4_4_in_pel.write = wr_line_buffer_3_4_out_pel.write;
        assign wr_fifo_mul_18_36_opA.write = wr_line_buffer_3_4_out_pel.write;     
        assign wr_fifo_line_buffer_4_5_in_pel.write = wr_line_buffer_3_5_out_pel.write;
        assign wr_fifo_mul_18_44_opA.write = wr_line_buffer_3_5_out_pel.write;
        assign wr_fifo_line_buffer_4_6_in_pel.write = wr_line_buffer_3_6_out_pel.write;
        assign wr_fifo_mul_18_52_opA.write = wr_line_buffer_3_6_out_pel.write;     
        assign wr_fifo_line_buffer_4_7_in_pel.write = wr_line_buffer_3_7_out_pel.write;
        assign wr_fifo_mul_18_60_opA.write = wr_line_buffer_3_7_out_pel.write;
                        
        // - DATA
        assign wr_fifo_line_buffer_4_0_in_pel.din = wr_line_buffer_3_0_out_pel.din;
        assign wr_fifo_mul_18_4_opA.din = wr_line_buffer_3_0_out_pel.din;
        assign wr_fifo_line_buffer_4_1_in_pel.din = wr_line_buffer_3_1_out_pel.din;
        assign wr_fifo_mul_18_12_opA.din = wr_line_buffer_3_1_out_pel.din;
        assign wr_fifo_line_buffer_4_2_in_pel.din = wr_line_buffer_3_2_out_pel.din;
        assign wr_fifo_mul_18_20_opA.din = wr_line_buffer_3_2_out_pel.din;     
        assign wr_fifo_line_buffer_4_3_in_pel.din = wr_line_buffer_3_3_out_pel.din;
        assign wr_fifo_mul_18_28_opA.din = wr_line_buffer_3_3_out_pel.din;
        assign wr_fifo_line_buffer_4_4_in_pel.din = wr_line_buffer_3_4_out_pel.din;
        assign wr_fifo_mul_18_36_opA.din = wr_line_buffer_3_4_out_pel.din;     
        assign wr_fifo_line_buffer_4_5_in_pel.din = wr_line_buffer_3_5_out_pel.din;
        assign wr_fifo_mul_18_44_opA.din = wr_line_buffer_3_5_out_pel.din;
        assign wr_fifo_line_buffer_4_6_in_pel.din = wr_line_buffer_3_6_out_pel.din;
        assign wr_fifo_mul_18_52_opA.din = wr_line_buffer_3_6_out_pel.din;     
        assign wr_fifo_line_buffer_4_7_in_pel.din = wr_line_buffer_3_7_out_pel.din;
        assign wr_fifo_mul_18_60_opA.din = wr_line_buffer_3_7_out_pel.din;
    
    //FORK line_buffer_4 to mul_18_5 & mul_18_13 & mul_18_21 & mul_18_29 & mul_18_37 & mul_18_45 & mul_18_53 & mul_18_61  

        // - INTERFACES 
        write_interface #(18,FLUX) wr_fifo_line_buffer_5_0_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_5_1_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_5_2_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_5_3_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_5_4_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_5_5_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_5_6_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_5_7_in_pel(clk);
        
        write_interface #(18,FLUX) wr_fifo_mul_18_5_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_13_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_21_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_29_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_37_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_45_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_53_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_61_opA(clk);               
     
        // - FULL
        assign wr_line_buffer_4_0_out_pel.full = wr_fifo_line_buffer_5_0_in_pel.full | wr_fifo_mul_18_5_opA.full;
        assign wr_line_buffer_4_1_out_pel.full = wr_fifo_line_buffer_5_1_in_pel.full | wr_fifo_mul_18_13_opA.full;
        assign wr_line_buffer_4_2_out_pel.full = wr_fifo_line_buffer_5_2_in_pel.full | wr_fifo_mul_18_21_opA.full;
        assign wr_line_buffer_4_3_out_pel.full = wr_fifo_line_buffer_5_3_in_pel.full | wr_fifo_mul_18_29_opA.full;
        assign wr_line_buffer_4_4_out_pel.full = wr_fifo_line_buffer_5_4_in_pel.full | wr_fifo_mul_18_37_opA.full;
        assign wr_line_buffer_4_5_out_pel.full = wr_fifo_line_buffer_5_5_in_pel.full | wr_fifo_mul_18_45_opA.full;
        assign wr_line_buffer_4_6_out_pel.full = wr_fifo_line_buffer_5_6_in_pel.full | wr_fifo_mul_18_53_opA.full;
        assign wr_line_buffer_4_7_out_pel.full = wr_fifo_line_buffer_5_7_in_pel.full | wr_fifo_mul_18_61_opA.full;
     
        // - WRITE
        assign wr_fifo_line_buffer_5_0_in_pel.write = wr_line_buffer_4_0_out_pel.write;
        assign wr_fifo_mul_18_5_opA.write = wr_line_buffer_4_0_out_pel.write;
        assign wr_fifo_line_buffer_5_1_in_pel.write = wr_line_buffer_4_1_out_pel.write;
        assign wr_fifo_mul_18_13_opA.write = wr_line_buffer_4_1_out_pel.write;
        assign wr_fifo_line_buffer_5_2_in_pel.write = wr_line_buffer_4_2_out_pel.write;
        assign wr_fifo_mul_18_21_opA.write = wr_line_buffer_4_2_out_pel.write;     
        assign wr_fifo_line_buffer_5_3_in_pel.write = wr_line_buffer_4_3_out_pel.write;
        assign wr_fifo_mul_18_29_opA.write = wr_line_buffer_4_3_out_pel.write;
        assign wr_fifo_line_buffer_5_4_in_pel.write = wr_line_buffer_4_4_out_pel.write;
        assign wr_fifo_mul_18_37_opA.write = wr_line_buffer_4_4_out_pel.write;     
        assign wr_fifo_line_buffer_5_5_in_pel.write = wr_line_buffer_4_5_out_pel.write;
        assign wr_fifo_mul_18_45_opA.write = wr_line_buffer_4_5_out_pel.write;
        assign wr_fifo_line_buffer_5_6_in_pel.write = wr_line_buffer_4_6_out_pel.write;
        assign wr_fifo_mul_18_53_opA.write = wr_line_buffer_4_6_out_pel.write;     
        assign wr_fifo_line_buffer_5_7_in_pel.write = wr_line_buffer_4_7_out_pel.write;
        assign wr_fifo_mul_18_61_opA.write = wr_line_buffer_4_7_out_pel.write;
                        
        // - DATA
        assign wr_fifo_line_buffer_5_0_in_pel.din = wr_line_buffer_4_0_out_pel.din;
        assign wr_fifo_mul_18_5_opA.din = wr_line_buffer_4_0_out_pel.din;
        assign wr_fifo_line_buffer_5_1_in_pel.din = wr_line_buffer_4_1_out_pel.din;
        assign wr_fifo_mul_18_13_opA.din = wr_line_buffer_4_1_out_pel.din;
        assign wr_fifo_line_buffer_5_2_in_pel.din = wr_line_buffer_4_2_out_pel.din;
        assign wr_fifo_mul_18_21_opA.din = wr_line_buffer_4_2_out_pel.din;     
        assign wr_fifo_line_buffer_5_3_in_pel.din = wr_line_buffer_4_3_out_pel.din;
        assign wr_fifo_mul_18_29_opA.din = wr_line_buffer_4_3_out_pel.din;
        assign wr_fifo_line_buffer_5_4_in_pel.din = wr_line_buffer_4_4_out_pel.din;
        assign wr_fifo_mul_18_37_opA.din = wr_line_buffer_4_4_out_pel.din;     
        assign wr_fifo_line_buffer_5_5_in_pel.din = wr_line_buffer_4_5_out_pel.din;
        assign wr_fifo_mul_18_45_opA.din = wr_line_buffer_4_5_out_pel.din;
        assign wr_fifo_line_buffer_5_6_in_pel.din = wr_line_buffer_4_6_out_pel.din;
        assign wr_fifo_mul_18_53_opA.din = wr_line_buffer_4_6_out_pel.din;     
        assign wr_fifo_line_buffer_5_7_in_pel.din = wr_line_buffer_4_7_out_pel.din;
        assign wr_fifo_mul_18_61_opA.din = wr_line_buffer_4_7_out_pel.din;
        
    //FORK line_buffer_5 to mul_18_6 & mul_18_14 & mul_18_22 & mul_18_30 & mul_18_38 & mul_18_46 & mul_18_54 & mul_18_62

        // - INTERFACES 
        write_interface #(18,FLUX) wr_fifo_line_buffer_6_0_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_6_1_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_6_2_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_6_3_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_6_4_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_6_5_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_6_6_in_pel(clk);
        write_interface #(18,FLUX) wr_fifo_line_buffer_6_7_in_pel(clk);
        
        write_interface #(18,FLUX) wr_fifo_mul_18_6_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_14_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_22_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_30_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_38_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_46_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_54_opA(clk);
        write_interface #(18,FLUX) wr_fifo_mul_18_62_opA(clk);               
     
        // - FULL
        assign wr_line_buffer_5_0_out_pel.full = wr_fifo_line_buffer_6_0_in_pel.full | wr_fifo_mul_18_6_opA.full;
        assign wr_line_buffer_5_1_out_pel.full = wr_fifo_line_buffer_6_1_in_pel.full | wr_fifo_mul_18_14_opA.full;
        assign wr_line_buffer_5_2_out_pel.full = wr_fifo_line_buffer_6_2_in_pel.full | wr_fifo_mul_18_22_opA.full;
        assign wr_line_buffer_5_3_out_pel.full = wr_fifo_line_buffer_6_3_in_pel.full | wr_fifo_mul_18_30_opA.full;
        assign wr_line_buffer_5_4_out_pel.full = wr_fifo_line_buffer_6_4_in_pel.full | wr_fifo_mul_18_38_opA.full;
        assign wr_line_buffer_5_5_out_pel.full = wr_fifo_line_buffer_6_5_in_pel.full | wr_fifo_mul_18_46_opA.full;
        assign wr_line_buffer_5_6_out_pel.full = wr_fifo_line_buffer_6_6_in_pel.full | wr_fifo_mul_18_54_opA.full;
        assign wr_line_buffer_5_7_out_pel.full = wr_fifo_line_buffer_6_7_in_pel.full | wr_fifo_mul_18_62_opA.full;
     
        // - WRITE
        assign wr_fifo_line_buffer_6_0_in_pel.write = wr_line_buffer_5_0_out_pel.write;
        assign wr_fifo_mul_18_6_opA.write = wr_line_buffer_5_0_out_pel.write;
        assign wr_fifo_line_buffer_6_1_in_pel.write = wr_line_buffer_5_1_out_pel.write;
        assign wr_fifo_mul_18_14_opA.write = wr_line_buffer_5_1_out_pel.write;
        assign wr_fifo_line_buffer_6_2_in_pel.write = wr_line_buffer_5_2_out_pel.write;
        assign wr_fifo_mul_18_22_opA.write = wr_line_buffer_5_2_out_pel.write;     
        assign wr_fifo_line_buffer_6_3_in_pel.write = wr_line_buffer_5_3_out_pel.write;
        assign wr_fifo_mul_18_30_opA.write = wr_line_buffer_5_3_out_pel.write;
        assign wr_fifo_line_buffer_6_4_in_pel.write = wr_line_buffer_5_4_out_pel.write;
        assign wr_fifo_mul_18_38_opA.write = wr_line_buffer_5_4_out_pel.write;     
        assign wr_fifo_line_buffer_6_5_in_pel.write = wr_line_buffer_5_5_out_pel.write;
        assign wr_fifo_mul_18_46_opA.write = wr_line_buffer_5_5_out_pel.write;
        assign wr_fifo_line_buffer_6_6_in_pel.write = wr_line_buffer_5_6_out_pel.write;
        assign wr_fifo_mul_18_54_opA.write = wr_line_buffer_5_6_out_pel.write;     
        assign wr_fifo_line_buffer_6_7_in_pel.write = wr_line_buffer_5_7_out_pel.write;
        assign wr_fifo_mul_18_62_opA.write = wr_line_buffer_5_7_out_pel.write;
                        
        // - DATA
        assign wr_fifo_line_buffer_6_0_in_pel.din = wr_line_buffer_5_0_out_pel.din;
        assign wr_fifo_mul_18_6_opA.din = wr_line_buffer_5_0_out_pel.din;
        assign wr_fifo_line_buffer_6_1_in_pel.din = wr_line_buffer_5_1_out_pel.din;
        assign wr_fifo_mul_18_14_opA.din = wr_line_buffer_5_1_out_pel.din;
        assign wr_fifo_line_buffer_6_2_in_pel.din = wr_line_buffer_5_2_out_pel.din;
        assign wr_fifo_mul_18_22_opA.din = wr_line_buffer_5_2_out_pel.din;     
        assign wr_fifo_line_buffer_6_3_in_pel.din = wr_line_buffer_5_3_out_pel.din;
        assign wr_fifo_mul_18_30_opA.din = wr_line_buffer_5_3_out_pel.din;
        assign wr_fifo_line_buffer_6_4_in_pel.din = wr_line_buffer_5_4_out_pel.din;
        assign wr_fifo_mul_18_38_opA.din = wr_line_buffer_5_4_out_pel.din;     
        assign wr_fifo_line_buffer_6_5_in_pel.din = wr_line_buffer_5_5_out_pel.din;
        assign wr_fifo_mul_18_46_opA.din = wr_line_buffer_5_5_out_pel.din;
        assign wr_fifo_line_buffer_6_6_in_pel.din = wr_line_buffer_5_6_out_pel.din;
        assign wr_fifo_mul_18_54_opA.din = wr_line_buffer_5_6_out_pel.din;     
        assign wr_fifo_line_buffer_6_7_in_pel.din = wr_line_buffer_5_7_out_pel.din;
        assign wr_fifo_mul_18_62_opA.din = wr_line_buffer_5_7_out_pel.din;

    //FORK coeff v C0 TO mul_18_0 & mul_18_8 & mul_18_16 & MUL_24 & MUL_32 & MUL_40 & MUL_48 & MUL_56
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_18_0_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_8_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_18_16_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_24_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_32_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_40_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_48_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_56_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_v_c0.full = wr_fifo_mul_18_0_opB.full | wr_fifo_mul_18_8_opB.full | wr_fifo_mul_18_16_opB.full 
        | wr_fifo_mul_18_24_opB.full | wr_fifo_mul_18_32_opB.full | wr_fifo_mul_18_40_opB.full | wr_fifo_mul_18_48_opB.full
        | wr_fifo_mul_18_56_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_18_0_opB.write = wr_coeff_luma_v_c0.write;
        assign wr_fifo_mul_18_8_opB.write = wr_coeff_luma_v_c0.write;
        assign wr_fifo_mul_18_16_opB.write = wr_coeff_luma_v_c0.write;
        assign wr_fifo_mul_18_24_opB.write = wr_coeff_luma_v_c0.write;
        assign wr_fifo_mul_18_32_opB.write = wr_coeff_luma_v_c0.write;
        assign wr_fifo_mul_18_40_opB.write = wr_coeff_luma_v_c0.write;
        assign wr_fifo_mul_18_48_opB.write = wr_coeff_luma_v_c0.write;
        assign wr_fifo_mul_18_56_opB.write = wr_coeff_luma_v_c0.write;
        
        // - DATA
        assign wr_fifo_mul_18_0_opB.din = wr_coeff_luma_v_c0.din;
        assign wr_fifo_mul_18_8_opB.din = wr_coeff_luma_v_c0.din;
        assign wr_fifo_mul_18_16_opB.din = wr_coeff_luma_v_c0.din;
        assign wr_fifo_mul_18_24_opB.din = wr_coeff_luma_v_c0.din;
        assign wr_fifo_mul_18_32_opB.din = wr_coeff_luma_v_c0.din;
        assign wr_fifo_mul_18_40_opB.din = wr_coeff_luma_v_c0.din;
        assign wr_fifo_mul_18_48_opB.din = wr_coeff_luma_v_c0.din;
        assign wr_fifo_mul_18_56_opB.din = wr_coeff_luma_v_c0.din;
        
    //FORK coeff h C1 TO mul_18_1 & mul_18_9 & mul_18_17 & MUL_25 & MUL_33 & MUL_41 & MUL_49 & MUL_57
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_18_1_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_9_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_18_17_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_25_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_33_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_41_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_49_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_57_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_v_c1.full = wr_fifo_mul_18_1_opB.full | wr_fifo_mul_18_9_opB.full | wr_fifo_mul_18_17_opB.full 
        | wr_fifo_mul_18_25_opB.full | wr_fifo_mul_18_33_opB.full | wr_fifo_mul_18_41_opB.full | wr_fifo_mul_18_49_opB.full
        | wr_fifo_mul_18_57_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_18_1_opB.write = wr_coeff_luma_v_c1.write;
        assign wr_fifo_mul_18_9_opB.write = wr_coeff_luma_v_c1.write;
        assign wr_fifo_mul_18_17_opB.write = wr_coeff_luma_v_c1.write;
        assign wr_fifo_mul_18_25_opB.write = wr_coeff_luma_v_c1.write;
        assign wr_fifo_mul_18_33_opB.write = wr_coeff_luma_v_c1.write;
        assign wr_fifo_mul_18_41_opB.write = wr_coeff_luma_v_c1.write;
        assign wr_fifo_mul_18_49_opB.write = wr_coeff_luma_v_c1.write;
        assign wr_fifo_mul_18_57_opB.write = wr_coeff_luma_v_c1.write;
        
        // - DATA
        assign wr_fifo_mul_18_1_opB.din = wr_coeff_luma_v_c1.din;
        assign wr_fifo_mul_18_9_opB.din = wr_coeff_luma_v_c1.din;
        assign wr_fifo_mul_18_17_opB.din = wr_coeff_luma_v_c1.din;
        assign wr_fifo_mul_18_25_opB.din = wr_coeff_luma_v_c1.din;
        assign wr_fifo_mul_18_33_opB.din = wr_coeff_luma_v_c1.din;
        assign wr_fifo_mul_18_41_opB.din = wr_coeff_luma_v_c1.din;
        assign wr_fifo_mul_18_49_opB.din = wr_coeff_luma_v_c1.din;
        assign wr_fifo_mul_18_57_opB.din = wr_coeff_luma_v_c1.din;            
    
    //FORK coeff h C2 TO mul_18_2 & mul_18_10 & mul_18_18 & MUL_26 & MUL_34 & MUL_42 & MUL_50 & MUL_58
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_18_2_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_10_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_18_18_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_26_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_34_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_42_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_50_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_58_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_v_c2.full = wr_fifo_mul_18_2_opB.full | wr_fifo_mul_18_10_opB.full | wr_fifo_mul_18_18_opB.full 
        | wr_fifo_mul_18_26_opB.full | wr_fifo_mul_18_34_opB.full | wr_fifo_mul_18_42_opB.full | wr_fifo_mul_18_50_opB.full
        | wr_fifo_mul_18_58_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_18_2_opB.write = wr_coeff_luma_v_c2.write;
        assign wr_fifo_mul_18_10_opB.write = wr_coeff_luma_v_c2.write;
        assign wr_fifo_mul_18_18_opB.write = wr_coeff_luma_v_c2.write;
        assign wr_fifo_mul_18_26_opB.write = wr_coeff_luma_v_c2.write;
        assign wr_fifo_mul_18_34_opB.write = wr_coeff_luma_v_c2.write;
        assign wr_fifo_mul_18_42_opB.write = wr_coeff_luma_v_c2.write;
        assign wr_fifo_mul_18_50_opB.write = wr_coeff_luma_v_c2.write;
        assign wr_fifo_mul_18_58_opB.write = wr_coeff_luma_v_c2.write;
        
        // - DATA
        assign wr_fifo_mul_18_2_opB.din = wr_coeff_luma_v_c2.din;
        assign wr_fifo_mul_18_10_opB.din = wr_coeff_luma_v_c2.din;
        assign wr_fifo_mul_18_18_opB.din = wr_coeff_luma_v_c2.din;
        assign wr_fifo_mul_18_26_opB.din = wr_coeff_luma_v_c2.din;
        assign wr_fifo_mul_18_34_opB.din = wr_coeff_luma_v_c2.din;
        assign wr_fifo_mul_18_42_opB.din = wr_coeff_luma_v_c2.din;
        assign wr_fifo_mul_18_50_opB.din = wr_coeff_luma_v_c2.din;
        assign wr_fifo_mul_18_58_opB.din = wr_coeff_luma_v_c2.din;
        
    //FORK coeff h C3 TO mul_18_3 & mul_18_11 & mul_18_19 & MUL_27 & MUL_35 & MUL_43 & MUL_51 & MUL_59
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_18_3_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_11_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_18_19_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_27_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_35_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_43_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_51_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_59_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_v_c3.full = wr_fifo_mul_18_3_opB.full | wr_fifo_mul_18_11_opB.full | wr_fifo_mul_18_19_opB.full 
        | wr_fifo_mul_18_27_opB.full | wr_fifo_mul_18_35_opB.full | wr_fifo_mul_18_43_opB.full | wr_fifo_mul_18_51_opB.full
        | wr_fifo_mul_18_59_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_18_3_opB.write = wr_coeff_luma_v_c3.write;
        assign wr_fifo_mul_18_11_opB.write = wr_coeff_luma_v_c3.write;
        assign wr_fifo_mul_18_19_opB.write = wr_coeff_luma_v_c3.write;
        assign wr_fifo_mul_18_27_opB.write = wr_coeff_luma_v_c3.write;
        assign wr_fifo_mul_18_35_opB.write = wr_coeff_luma_v_c3.write;
        assign wr_fifo_mul_18_43_opB.write = wr_coeff_luma_v_c3.write;
        assign wr_fifo_mul_18_51_opB.write = wr_coeff_luma_v_c3.write;
        assign wr_fifo_mul_18_59_opB.write = wr_coeff_luma_v_c3.write;
        
        // - DATA
        assign wr_fifo_mul_18_3_opB.din = wr_coeff_luma_v_c3.din;
        assign wr_fifo_mul_18_11_opB.din = wr_coeff_luma_v_c3.din;
        assign wr_fifo_mul_18_19_opB.din = wr_coeff_luma_v_c3.din;
        assign wr_fifo_mul_18_27_opB.din = wr_coeff_luma_v_c3.din;
        assign wr_fifo_mul_18_35_opB.din = wr_coeff_luma_v_c3.din;
        assign wr_fifo_mul_18_43_opB.din = wr_coeff_luma_v_c3.din;
        assign wr_fifo_mul_18_51_opB.din = wr_coeff_luma_v_c3.din;
        assign wr_fifo_mul_18_59_opB.din = wr_coeff_luma_v_c3.din;        

    //FORK coeff h C4 TO mul_18_4 & mul_18_12 & mul_18_20 & MUL_28 & MUL_36 & MUL_44 & MUL_52 & MUL_60
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_18_4_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_12_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_18_20_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_28_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_36_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_44_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_52_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_60_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_v_c4.full = wr_fifo_mul_18_4_opB.full | wr_fifo_mul_18_12_opB.full | wr_fifo_mul_18_20_opB.full 
        | wr_fifo_mul_18_28_opB.full | wr_fifo_mul_18_36_opB.full | wr_fifo_mul_18_44_opB.full | wr_fifo_mul_18_52_opB.full
        | wr_fifo_mul_18_60_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_18_4_opB.write = wr_coeff_luma_v_c4.write;
        assign wr_fifo_mul_18_12_opB.write = wr_coeff_luma_v_c4.write;
        assign wr_fifo_mul_18_20_opB.write = wr_coeff_luma_v_c4.write;
        assign wr_fifo_mul_18_28_opB.write = wr_coeff_luma_v_c4.write;
        assign wr_fifo_mul_18_36_opB.write = wr_coeff_luma_v_c4.write;
        assign wr_fifo_mul_18_44_opB.write = wr_coeff_luma_v_c4.write;
        assign wr_fifo_mul_18_52_opB.write = wr_coeff_luma_v_c4.write;
        assign wr_fifo_mul_18_60_opB.write = wr_coeff_luma_v_c4.write;
        
        // - DATA
        assign wr_fifo_mul_18_4_opB.din = wr_coeff_luma_v_c4.din;
        assign wr_fifo_mul_18_12_opB.din = wr_coeff_luma_v_c4.din;
        assign wr_fifo_mul_18_20_opB.din = wr_coeff_luma_v_c4.din;
        assign wr_fifo_mul_18_28_opB.din = wr_coeff_luma_v_c4.din;
        assign wr_fifo_mul_18_36_opB.din = wr_coeff_luma_v_c4.din;
        assign wr_fifo_mul_18_44_opB.din = wr_coeff_luma_v_c4.din;
        assign wr_fifo_mul_18_52_opB.din = wr_coeff_luma_v_c4.din;
        assign wr_fifo_mul_18_60_opB.din = wr_coeff_luma_v_c4.din;

    //FORK coeff h C5 TO mul_18_5 & mul_18_13 & mul_18_21 & MUL_29 & MUL_37 & MUL_45 & MUL_53 & MUL_61
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_18_5_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_13_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_18_21_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_29_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_37_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_45_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_53_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_61_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_v_c5.full = wr_fifo_mul_18_5_opB.full | wr_fifo_mul_18_13_opB.full | wr_fifo_mul_18_21_opB.full 
        | wr_fifo_mul_18_29_opB.full | wr_fifo_mul_18_37_opB.full | wr_fifo_mul_18_45_opB.full | wr_fifo_mul_18_53_opB.full
        | wr_fifo_mul_18_61_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_18_5_opB.write = wr_coeff_luma_v_c5.write;
        assign wr_fifo_mul_18_13_opB.write = wr_coeff_luma_v_c5.write;
        assign wr_fifo_mul_18_21_opB.write = wr_coeff_luma_v_c5.write;
        assign wr_fifo_mul_18_29_opB.write = wr_coeff_luma_v_c5.write;
        assign wr_fifo_mul_18_37_opB.write = wr_coeff_luma_v_c5.write;
        assign wr_fifo_mul_18_45_opB.write = wr_coeff_luma_v_c5.write;
        assign wr_fifo_mul_18_53_opB.write = wr_coeff_luma_v_c5.write;
        assign wr_fifo_mul_18_61_opB.write = wr_coeff_luma_v_c5.write;
        
        // - DATA
        assign wr_fifo_mul_18_5_opB.din = wr_coeff_luma_v_c5.din;
        assign wr_fifo_mul_18_13_opB.din = wr_coeff_luma_v_c5.din;
        assign wr_fifo_mul_18_21_opB.din = wr_coeff_luma_v_c5.din;
        assign wr_fifo_mul_18_29_opB.din = wr_coeff_luma_v_c5.din;
        assign wr_fifo_mul_18_37_opB.din = wr_coeff_luma_v_c5.din;
        assign wr_fifo_mul_18_45_opB.din = wr_coeff_luma_v_c5.din;
        assign wr_fifo_mul_18_53_opB.din = wr_coeff_luma_v_c5.din;
        assign wr_fifo_mul_18_61_opB.din = wr_coeff_luma_v_c5.din;
        
    //FORK coeff h C6 TO mul_18_6 & mul_18_14 & mul_18_22 & MUL_30 & MUL_38 & MUL_46 & MUL_54 & MUL_62
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_18_6_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_14_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_18_22_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_30_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_38_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_46_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_54_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_62_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_v_c6.full = wr_fifo_mul_18_6_opB.full | wr_fifo_mul_18_14_opB.full | wr_fifo_mul_18_22_opB.full 
        | wr_fifo_mul_18_30_opB.full | wr_fifo_mul_18_38_opB.full | wr_fifo_mul_18_46_opB.full | wr_fifo_mul_18_54_opB.full
        | wr_fifo_mul_18_62_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_18_6_opB.write = wr_coeff_luma_v_c6.write;
        assign wr_fifo_mul_18_14_opB.write = wr_coeff_luma_v_c6.write;
        assign wr_fifo_mul_18_22_opB.write = wr_coeff_luma_v_c6.write;
        assign wr_fifo_mul_18_30_opB.write = wr_coeff_luma_v_c6.write;
        assign wr_fifo_mul_18_38_opB.write = wr_coeff_luma_v_c6.write;
        assign wr_fifo_mul_18_46_opB.write = wr_coeff_luma_v_c6.write;
        assign wr_fifo_mul_18_54_opB.write = wr_coeff_luma_v_c6.write;
        assign wr_fifo_mul_18_62_opB.write = wr_coeff_luma_v_c6.write;
        
        // - DATA
        assign wr_fifo_mul_18_6_opB.din = wr_coeff_luma_v_c6.din;
        assign wr_fifo_mul_18_14_opB.din = wr_coeff_luma_v_c6.din;
        assign wr_fifo_mul_18_22_opB.din = wr_coeff_luma_v_c6.din;
        assign wr_fifo_mul_18_30_opB.din = wr_coeff_luma_v_c6.din;
        assign wr_fifo_mul_18_38_opB.din = wr_coeff_luma_v_c6.din;
        assign wr_fifo_mul_18_46_opB.din = wr_coeff_luma_v_c6.din;
        assign wr_fifo_mul_18_54_opB.din = wr_coeff_luma_v_c6.din;
        assign wr_fifo_mul_18_62_opB.din = wr_coeff_luma_v_c6.din;        

    //FORK coeff h C7 TO mul_18_7 & mul_18_15 & mul_18_23 & MUL_31 & MUL_39 & MUL_47 & MUL_55 & MUL_63
    
        // - INTERFACES   		    		
        write_interface #(9,FLUX) wr_fifo_mul_18_7_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_15_opB(clk); 
        write_interface #(9,FLUX) wr_fifo_mul_18_23_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_31_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_39_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_47_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_55_opB(clk);
        write_interface #(9,FLUX) wr_fifo_mul_18_63_opB(clk);                
                       
        // - FULL
        assign wr_coeff_luma_v_c7.full = wr_fifo_mul_18_7_opB.full | wr_fifo_mul_18_15_opB.full | wr_fifo_mul_18_23_opB.full 
        | wr_fifo_mul_18_31_opB.full | wr_fifo_mul_18_39_opB.full | wr_fifo_mul_18_47_opB.full | wr_fifo_mul_18_55_opB.full
        | wr_fifo_mul_18_63_opB.full;
        
        // - WRITE
        assign wr_fifo_mul_18_7_opB.write = wr_coeff_luma_v_c7.write;
        assign wr_fifo_mul_18_15_opB.write = wr_coeff_luma_v_c7.write;
        assign wr_fifo_mul_18_23_opB.write = wr_coeff_luma_v_c7.write;
        assign wr_fifo_mul_18_31_opB.write = wr_coeff_luma_v_c7.write;
        assign wr_fifo_mul_18_39_opB.write = wr_coeff_luma_v_c7.write;
        assign wr_fifo_mul_18_47_opB.write = wr_coeff_luma_v_c7.write;
        assign wr_fifo_mul_18_55_opB.write = wr_coeff_luma_v_c7.write;
        assign wr_fifo_mul_18_63_opB.write = wr_coeff_luma_v_c7.write;
        
        // - DATA
        assign wr_fifo_mul_18_7_opB.din = wr_coeff_luma_v_c7.din;
        assign wr_fifo_mul_18_15_opB.din = wr_coeff_luma_v_c7.din;
        assign wr_fifo_mul_18_23_opB.din = wr_coeff_luma_v_c7.din;
        assign wr_fifo_mul_18_31_opB.din = wr_coeff_luma_v_c7.din;
        assign wr_fifo_mul_18_39_opB.din = wr_coeff_luma_v_c7.din;
        assign wr_fifo_mul_18_47_opB.din = wr_coeff_luma_v_c7.din;
        assign wr_fifo_mul_18_55_opB.din = wr_coeff_luma_v_c7.din;
        assign wr_fifo_mul_18_63_opB.din = wr_coeff_luma_v_c7.din;



//FINE FORKS



    
//FIFO PRIMA PARTE 



    //extsize<->derive_real_size
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_derive_real_size
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_derive_real_size_ext_size.fifo),
        .read_port(rd_derive_real_size_ext_size.fifo)
        );
      
    //extsize<->remove_h_0
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_h_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_h_0_ext_size.fifo),
        .read_port(rd_remove_h_0_ext_size.fifo)
        );
		
	//extsize<->remove_h_1
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_h_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_h_1_ext_size.fifo),
        .read_port(rd_remove_h_1_ext_size.fifo)
        );
		
	//extsize<->remove_h_2
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_h_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_h_2_ext_size.fifo),
        .read_port(rd_remove_h_2_ext_size.fifo)
        );
		
	//extsize<->remove_h_3
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_h_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_h_3_ext_size.fifo),
        .read_port(rd_remove_h_3_ext_size.fifo)
        );
		
	//extsize<->remove_h_4
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_h_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_h_4_ext_size.fifo),
        .read_port(rd_remove_h_4_ext_size.fifo)
        );
		
	//extsize<->remove_h_5
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_h_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_h_5_ext_size.fifo),
        .read_port(rd_remove_h_5_ext_size.fifo)
        );
		
	//extsize<->remove_h_6
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_h_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_h_6_ext_size.fifo),
        .read_port(rd_remove_h_6_ext_size.fifo)
        );
		
	//extsize<->remove_h_7
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_h_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_h_7_ext_size.fifo),
        .read_port(rd_remove_h_7_ext_size.fifo)
        );
	
    
    //h_alpha<->coeff_h
        
        //h_alpha<->coeff_luma_h
        fifo_ms #(3,DEPTH,FLUX) fifo_h_alpha_coeff_luma_h_alpha
        (
        .clk(clk),
        .rst(rst),
        .write_port(write_port_h_alpha),
        .read_port(rd_coeff_luma_h_alpha.fifo)
        ); 
            
    //v_alpha<->coeff_v
    
        //v_aplha<->coeff_luma_v
        fifo_ms #(3,DEPTH,FLUX) fifo_v_alpha_coeff_luma_v_alpha
        (
        .clk(clk),
        .rst(rst),
        .write_port(write_port_v_alpha),
        .read_port(rd_coeff_luma_v_alpha.fifo)
        );


    //extsize mul9

    //1� riga                 
        //extsize<->mul_9_0        
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_0_ext_size.fifo),
        .read_port(rd_mul_9_0_ext_size.fifo)
        );        
                
        //extsize<->mul_9_1
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_1_ext_size.fifo),
        .read_port(rd_mul_9_1_ext_size.fifo)
        );
                
        //extsize<->mul_9_2
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_2_ext_size.fifo),
        .read_port(rd_mul_9_2_ext_size.fifo)
        );
        
        //extsize<->mul_9_3
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_3_ext_size.fifo),
        .read_port(rd_mul_9_3_ext_size.fifo)
        );
                
        //extsize<->mul_9_4
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_4_ext_size.fifo),
        .read_port(rd_mul_9_4_ext_size.fifo)
        );
        
        //extsize<->mul_9_5
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_5_ext_size.fifo),
        .read_port(rd_mul_9_5_ext_size.fifo)
        );        
        
        //extsize<->mul_9_6
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_6_ext_size.fifo),
        .read_port(rd_mul_9_6_ext_size.fifo)
        );
                
        //extsize<->mul_9_7
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_7_ext_size.fifo),
        .read_port(rd_mul_9_7_ext_size.fifo)
        );
  
    //2�riga
                   
        //extsize<->mul_9_8        
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_8
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_8_ext_size.fifo),
        .read_port(rd_mul_9_8_ext_size.fifo)
        );        
                
        //extsize<->mul_9_9
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_9
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_9_ext_size.fifo),
        .read_port(rd_mul_9_9_ext_size.fifo)
        );
                
        //extsize<->mul_9_10
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_10
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_10_ext_size.fifo),
        .read_port(rd_mul_9_10_ext_size.fifo)
        );
        
        //extsize<->mul_9_11
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_11
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_11_ext_size.fifo),
        .read_port(rd_mul_9_11_ext_size.fifo)
        );
                
        //extsize<->mul_9_12
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_12
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_12_ext_size.fifo),
        .read_port(rd_mul_9_12_ext_size.fifo)
        );
        
        //extsize<->mul_9_13
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_13
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_13_ext_size.fifo),
        .read_port(rd_mul_9_13_ext_size.fifo)
        );        
        
        //extsize<->mul_9_14
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_14
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_14_ext_size.fifo),
        .read_port(rd_mul_9_14_ext_size.fifo)
        );
                
        //extsize<->mul_9_15
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_15
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_15_ext_size.fifo),
        .read_port(rd_mul_9_15_ext_size.fifo)
        );
  
    //3�riga
                 
        //extsize<->mul_9_16        
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_16
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_16_ext_size.fifo),
        .read_port(rd_mul_9_16_ext_size.fifo)
        );        
                
        //extsize<->mul_9_17
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_17
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_17_ext_size.fifo),
        .read_port(rd_mul_9_17_ext_size.fifo)
        );
                
        //extsize<->mul_9_18
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_18
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_18_ext_size.fifo),
        .read_port(rd_mul_9_18_ext_size.fifo)
        );
        
        //extsize<->mul_9_19
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_19
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_19_ext_size.fifo),
        .read_port(rd_mul_9_19_ext_size.fifo)
        );
                
        //extsize<->mul_9_20
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_20
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_20_ext_size.fifo),
        .read_port(rd_mul_9_20_ext_size.fifo)
        );
        
        //extsize<->mul_9_21
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_21
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_21_ext_size.fifo),
        .read_port(rd_mul_9_21_ext_size.fifo)
        );        
        
        //extsize<->mul_9_22
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_22
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_22_ext_size.fifo),
        .read_port(rd_mul_9_22_ext_size.fifo)
        );
                
        //extsize<->mul_9_23
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_23
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_23_ext_size.fifo),
        .read_port(rd_mul_9_23_ext_size.fifo)
        );
    
    //4�riga
                     
        //extsize<->mul_9_24        
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_24
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_24_ext_size.fifo),
        .read_port(rd_mul_9_24_ext_size.fifo)
        );        
                
        //extsize<->mul_9_25
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_25
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_25_ext_size.fifo),
        .read_port(rd_mul_9_25_ext_size.fifo)
        );
                
        //extsize<->mul_9_26
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_26
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_26_ext_size.fifo),
        .read_port(rd_mul_9_26_ext_size.fifo)
        );
        
        //extsize<->mul_9_27
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_27
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_27_ext_size.fifo),
        .read_port(rd_mul_9_27_ext_size.fifo)
        );
                
        //extsize<->mul_9_28
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_28
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_28_ext_size.fifo),
        .read_port(rd_mul_9_28_ext_size.fifo)
        );
        
        //extsize<->mul_9_29
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_29
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_29_ext_size.fifo),
        .read_port(rd_mul_9_29_ext_size.fifo)
        );        
        
        //extsize<->mul_9_30
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_30
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_30_ext_size.fifo),
        .read_port(rd_mul_9_30_ext_size.fifo)
        );
                
        //extsize<->mul_9_31
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_31
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_31_ext_size.fifo),
        .read_port(rd_mul_9_31_ext_size.fifo)
        );
            
    //5�riga

        //extsize<->mul_9_32
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_32
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_32_ext_size.fifo),
        .read_port(rd_mul_9_32_ext_size.fifo)
        );        
                
        //extsize<->mul_9_33
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_33
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_33_ext_size.fifo),
        .read_port(rd_mul_9_33_ext_size.fifo)
        );
                
        //extsize<->mul_9_34
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_34
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_34_ext_size.fifo),
        .read_port(rd_mul_9_34_ext_size.fifo)
        );
        
        //extsize<->mul_9_35
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_35
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_35_ext_size.fifo),
        .read_port(rd_mul_9_35_ext_size.fifo)
        );
                
        //extsize<->mul_9_36
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_36
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_36_ext_size.fifo),
        .read_port(rd_mul_9_36_ext_size.fifo)
        );
        
        //extsize<->mul_9_37
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_37
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_37_ext_size.fifo),
        .read_port(rd_mul_9_37_ext_size.fifo)
        );        
        
        //extsize<->mul_9_38
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_38
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_38_ext_size.fifo),
        .read_port(rd_mul_9_38_ext_size.fifo)
        );
                
        //extsize<->mul_9_39
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_39
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_39_ext_size.fifo),
        .read_port(rd_mul_9_39_ext_size.fifo)
        );
    
    //6�riga
        
        //extsize<->mul_9_40
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_40
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_40_ext_size.fifo),
        .read_port(rd_mul_9_40_ext_size.fifo)
        );        
                
        //extsize<->mul_9_41
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_41
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_41_ext_size.fifo),
        .read_port(rd_mul_9_41_ext_size.fifo)
        );
                
        //extsize<->mul_9_42
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_42
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_42_ext_size.fifo),
        .read_port(rd_mul_9_42_ext_size.fifo)
        );
        
        //extsize<->mul_9_43
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_43
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_43_ext_size.fifo),
        .read_port(rd_mul_9_43_ext_size.fifo)
        );
                
        //extsize<->mul_9_44
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_44
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_44_ext_size.fifo),
        .read_port(rd_mul_9_44_ext_size.fifo)
        );
        
        //extsize<->mul_9_45
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_45
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_45_ext_size.fifo),
        .read_port(rd_mul_9_45_ext_size.fifo)
        );        
        
        //extsize<->mul_9_46
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_46
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_46_ext_size.fifo),
        .read_port(rd_mul_9_46_ext_size.fifo)
        );
                
        //extsize<->mul_9_47
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_47
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_47_ext_size.fifo),
        .read_port(rd_mul_9_47_ext_size.fifo)
        );
    
    //7�riga
        
        //extsize<->mul_9_48
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_48
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_48_ext_size.fifo),
        .read_port(rd_mul_9_48_ext_size.fifo)
        );        
                
        //extsize<->mul_9_49
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_49
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_49_ext_size.fifo),
        .read_port(rd_mul_9_49_ext_size.fifo)
        );
                
        //extsize<->mul_9_50
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_50
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_50_ext_size.fifo),
        .read_port(rd_mul_9_50_ext_size.fifo)
        );
        
        //extsize<->mul_9_51
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_51
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_51_ext_size.fifo),
        .read_port(rd_mul_9_51_ext_size.fifo)
        );
                
        //extsize<->mul_9_52
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_52
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_52_ext_size.fifo),
        .read_port(rd_mul_9_52_ext_size.fifo)
        );
        
        //extsize<->mul_9_53
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_53
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_53_ext_size.fifo),
        .read_port(rd_mul_9_53_ext_size.fifo)
        );        
        
        //extsize<->mul_9_54
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_54
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_54_ext_size.fifo),
        .read_port(rd_mul_9_54_ext_size.fifo)
        );
                
        //extsize<->mul_9_55
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_55
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_55_ext_size.fifo),
        .read_port(rd_mul_9_55_ext_size.fifo)
        );    
    
    //8�riga
        
        //extsize<->mul_9_56
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_56
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_56_ext_size.fifo),
        .read_port(rd_mul_9_56_ext_size.fifo)
        );        
                
        //extsize<->mul_9_57
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_57
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_57_ext_size.fifo),
        .read_port(rd_mul_9_57_ext_size.fifo)
        );
                
        //extsize<->mul_9_58
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_58
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_58_ext_size.fifo),
        .read_port(rd_mul_9_58_ext_size.fifo)
        );
        
        //extsize<->mul_9_59
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_59
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_59_ext_size.fifo),
        .read_port(rd_mul_9_59_ext_size.fifo)
        );
                
        //extsize<->mul_9_60
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_60
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_60_ext_size.fifo),
        .read_port(rd_mul_9_60_ext_size.fifo)
        );
        
        //extsize<->mul_9_61
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_61
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_61_ext_size.fifo),
        .read_port(rd_mul_9_61_ext_size.fifo)
        );        
        
        //extsize<->mul_9_62
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_62
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_62_ext_size.fifo),
        .read_port(rd_mul_9_62_ext_size.fifo)
        );
                
        //extsize<->mul_9_63
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul9_63
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_63_ext_size.fifo),
        .read_port(rd_mul_9_63_ext_size.fifo)
        );

    //Blocco rosso fifo nel ppt
   
        //in_port_1<->delay_0
        fifo_ms #(8,DEPTH,FLUX) fifo_in_port_1_delay_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_delay_0_in_pel.fifo),
        .read_port(rd_delay_0_in_pel.fifo)
        );
		
        //in_port_2<->delay_1
        fifo_ms #(8,DEPTH,FLUX) fifo_in_port_2_delay_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_delay_1_in_pel.fifo),
        .read_port(rd_delay_1_in_pel.fifo)
        );

        //in_port_3<->delay_2
        fifo_ms #(8,DEPTH,FLUX) fifo_in_port_3_delay_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_delay_2_in_pel.fifo),
        .read_port(rd_delay_2_in_pel.fifo)
        );

        //in_port_4<->delay_3
        fifo_ms #(8,DEPTH,FLUX) fifo_in_port_4_delay_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_delay_3_in_pel.fifo),
        .read_port(rd_delay_3_in_pel.fifo)
        );

        //in_port_5<->delay_4
        fifo_ms #(8,DEPTH,FLUX) fifo_in_port_5_delay_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_delay_4_in_pel.fifo),
        .read_port(rd_delay_4_in_pel.fifo)
        );
		
        //in_port_6<->delay_5
        fifo_ms #(8,DEPTH,FLUX) fifo_in_port_6_delay_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_delay_5_in_pel.fifo),
        .read_port(rd_delay_5_in_pel.fifo)
        );		
		
        //in_port_7<->delay_6
        fifo_ms #(8,DEPTH,FLUX) fifo_in_port_7_delay_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_delay_6_in_pel.fifo),
        .read_port(rd_delay_6_in_pel.fifo)
        );		   
   
	//FIFO OPA <-> MUL_9_0 

	//input 0

        //inport0<->mul_9_0
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_0_mul_9_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_0_opA.fifo), 
        .read_port(rd_mul_9_0_opA.fifo)
        );

        //inport0<->mul9_15
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_0_mul_9_15
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_15_opA.fifo),
        .read_port(rd_mul_9_15_opA.fifo)
        );        
        
        //inport0<->mul9_22
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_0_mul_9_22
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_22_opA.fifo),
        .read_port(rd_mul_9_22_opA.fifo)
        );
        
        //inport0<->mul9_29
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_0_mul_9_29
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_29_opA.fifo),
        .read_port(rd_mul_9_29_opA.fifo)
        );

        //inport0<->mul9_36
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_0_mul_9_36
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_36_opA.fifo),
        .read_port(rd_mul_9_36_opA.fifo)
        );

        //inport0<->mul9_43
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_0_mul_9_43
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_43_opA.fifo),
        .read_port(rd_mul_9_43_opA.fifo)
        );

        //inport0<->mul9_50
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_0_mul_9_50
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_50_opA.fifo),
        .read_port(rd_mul_9_50_opA.fifo)
        );

        //inport0<->mul9_57
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_0_mul_9_57
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_57_opA.fifo),
        .read_port(rd_mul_9_57_opA.fifo)
        );    

	
	//input 1

        //inport1<->mul9_1
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_1_mul_9_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_1_opA.fifo),
        .read_port(rd_mul_9_1_opA.fifo)
        );
		                          
        //inport1<->mul9_23
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_1_mul_9_23
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_23_opA.fifo),
        .read_port(rd_mul_9_23_opA.fifo)
        );
        
        //inport1<->mul9_30
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_1_mul_9_30
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_30_opA.fifo),
        .read_port(rd_mul_9_30_opA.fifo)
        );

        //inport1<->mul9_37
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_1_mul_9_37
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_37_opA.fifo),
        .read_port(rd_mul_9_37_opA.fifo)
        );

        //inport1<->mul9_44
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_1_mul_9_44
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_44_opA.fifo),
        .read_port(rd_mul_9_44_opA.fifo)
        );

        //inport1<->mul9_51
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_1_mul_9_51
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_51_opA.fifo),
        .read_port(rd_mul_9_51_opA.fifo)
        );

        //inport1<->mul9_58
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_1_mul_9_58
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_58_opA.fifo),
        .read_port(rd_mul_9_58_opA.fifo)
        );		
	
	//input 2

        //inport2<->mul9_2
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_2_mul_9_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_2_opA.fifo),
        .read_port(rd_mul_9_2_opA.fifo)
        );

        //inport2<->mul9_31
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_2_mul_9_31
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_31_opA.fifo),
        .read_port(rd_mul_9_31_opA.fifo)
        );

        //inport2<->mul9_38
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_2_mul_9_38
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_38_opA.fifo),
        .read_port(rd_mul_9_38_opA.fifo)
        );

        //inport2<->mul9_45
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_2_mul_9_45
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_45_opA.fifo),
        .read_port(rd_mul_9_45_opA.fifo)
        );

        //inport2<->mul9_52
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_2_mul_9_52
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_52_opA.fifo),
        .read_port(rd_mul_9_52_opA.fifo)
        );

        //inport2<->mul9_59
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_2_mul_9_59
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_59_opA.fifo),
        .read_port(rd_mul_9_59_opA.fifo)
        );
	
	//input 3

        //inport3<->mul9_3
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_3_mul_9_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_3_opA.fifo),
        .read_port(rd_mul_9_3_opA.fifo)
        );

        //inport3<->mul9_39
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_3_mul_9_39
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_39_opA.fifo),
        .read_port(rd_mul_9_39_opA.fifo)
        );

        //inport3<->mul9_46
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_3_mul_9_46
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_46_opA.fifo),
        .read_port(rd_mul_9_46_opA.fifo)
        );

        //inport3<->mul9_53
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_3_mul_9_53
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_53_opA.fifo),
        .read_port(rd_mul_9_53_opA.fifo)
        );

        //inport3<->mul9_60
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_3_mul_9_60
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_60_opA.fifo),
        .read_port(rd_mul_9_60_opA.fifo)
        );
	
	//input 4

        //inport4<->mul9_4
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_4_mul_9_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_4_opA.fifo),
        .read_port(rd_mul_9_4_opA.fifo)
        );

        //inport4<->mul9_47
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_4_mul_9_47
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_47_opA.fifo),
        .read_port(rd_mul_9_47_opA.fifo)
        );

        //inport4<->mul9_54
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_4_mul_9_54
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_54_opA.fifo),
        .read_port(rd_mul_9_54_opA.fifo)
        );

        //inport4<->mul9_61
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_4_mul_9_61
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_61_opA.fifo),
        .read_port(rd_mul_9_61_opA.fifo)
        );
	
	//input 5

        //inport5<->mul9_5
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_5_mul_9_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_5_opA.fifo),
        .read_port(rd_mul_9_5_opA.fifo)
        );
	
        //inport5<->mul9_55
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_5_mul_9_55
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_55_opA.fifo),
        .read_port(rd_mul_9_55_opA.fifo)
        );

        //inport5<->mul9_62
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_5_mul_9_62
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_62_opA.fifo),
        .read_port(rd_mul_9_62_opA.fifo)
        );
	
	//input 6

        //inport6<->mul9_6
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_6_mul_9_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_6_opA.fifo),
        .read_port(rd_mul_9_6_opA.fifo)
        );

        //inport6<->mul9_63
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_6_mul_9_63
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_63_opA.fifo), 
        .read_port(rd_mul_9_63_opA.fifo)
        );
	
	//input 7 

        //inport7<->mul9_7
        fifo_ms #(8,DEPTH,FLUX) fifo_inport_7_mul_9_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_7_opA.fifo),
        .read_port(rd_mul_9_7_opA.fifo)
        );
	
	//delay0  (NO FORK)
	
        //delay0<->mul9_8
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_0_mul_9_8
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_delay_0_out_pel.fifo),
        .read_port(rd_mul_9_8_opA.fifo)
        );	
	
	//delay1

        //delay1<->mul9_9
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_1_mul_9_9
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_9_opA.fifo),
        .read_port(rd_mul_9_9_opA.fifo)
        );

        //delay1<->mul9_16
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_1_mul_9_16
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_16_opA.fifo),
        .read_port(rd_mul_9_16_opA.fifo)
        );
	
	//delay2

        //delay2<->mul9_10
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_2_mul_9_10
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_10_opA.fifo),
        .read_port(rd_mul_9_10_opA.fifo)
        );

        //delay2<->mul9_17
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_2_mul_9_17
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_17_opA.fifo),
        .read_port(rd_mul_9_17_opA.fifo)
        );
        
        //delay2<->mul9_24
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_2_mul_9_24
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_24_opA.fifo),
        .read_port(rd_mul_9_24_opA.fifo)
        );
	
	//delay3

        //delay3<->mul9_11
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_3_mul_9_11
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_11_opA.fifo),
        .read_port(rd_mul_9_11_opA.fifo)
        );        
        
        //delay3<->mul9_18
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_3_mul_9_18
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_18_opA.fifo),
        .read_port(rd_mul_9_18_opA.fifo)
        );
        
        //delay3<->mul9_25
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_3_mul_9_25
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_25_opA.fifo),
        .read_port(rd_mul_9_25_opA.fifo)
        );

        //delay3<->mul9_32
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_3_mul_9_32
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_32_opA.fifo),
        .read_port(rd_mul_9_32_opA.fifo)
        );
	
	//delay4

        //delay4<->mul9_12
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_4_mul_9_12
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_12_opA.fifo),
        .read_port(rd_mul_9_12_opA.fifo)
        );        
        
        //delay4<->mul9_19
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_4_mul_9_19
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_19_opA.fifo),
        .read_port(rd_mul_9_19_opA.fifo)
        );
        
        //delay4<->mul9_26
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_4_mul_9_26
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_26_opA.fifo),
        .read_port(rd_mul_9_26_opA.fifo)
        );

        //delay4<->mul9_33
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_4_mul_9_33
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_33_opA.fifo),
        .read_port(rd_mul_9_33_opA.fifo)
        );

        //delay4<->mul9_40
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_4_mul_9_40
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_40_opA.fifo),
        .read_port(rd_mul_9_40_opA.fifo)
        );
	
	//delay5

        //delay5<->mul9_13
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_5_mul_9_13
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_13_opA.fifo),
        .read_port(rd_mul_9_13_opA.fifo)
        );        
        
        //delay5<->mul9_20
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_5_mul_9_20
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_20_opA.fifo),
        .read_port(rd_mul_9_20_opA.fifo)
        );
        
        //delay5<->mul9_27
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_5_mul_9_27
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_27_opA.fifo),
        .read_port(rd_mul_9_27_opA.fifo)
        );

        //delay5<->mul9_34
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_5_mul_9_34
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_34_opA.fifo),
        .read_port(rd_mul_9_34_opA.fifo)
        );

        //delay5<->mul9_41
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_5_mul_9_41
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_41_opA.fifo),
        .read_port(rd_mul_9_41_opA.fifo)
        );

        //delay5<->mul9_48
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_5_mul_9_48
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_48_opA.fifo),
        .read_port(rd_mul_9_48_opA.fifo)
        );
	
	//delay6
	
        //delay6<->mul9_14
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_6_mul_9_14
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_14_opA.fifo),
        .read_port(rd_mul_9_14_opA.fifo)
        );        
        
        //delay6<->mul9_21
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_6_mul_9_21
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_21_opA.fifo),
        .read_port(rd_mul_9_21_opA.fifo)
        );
        
        //delay6<->mul9_28
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_6_mul_9_28
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_28_opA.fifo),
        .read_port(rd_mul_9_28_opA.fifo)
        );

        //delay6<->mul9_35
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_6_mul_9_35
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_35_opA.fifo),
        .read_port(rd_mul_9_35_opA.fifo)
        );

        //delay6<->mul9_42
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_6_mul_9_42
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_42_opA.fifo),
        .read_port(rd_mul_9_42_opA.fifo)
        );

        //delay6<->mul9_49
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_6_mul_9_49
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_49_opA.fifo),
        .read_port(rd_mul_9_49_opA.fifo)
        );

        //delay6<->mul9_56
        fifo_ms #(8,DEPTH,FLUX) fifo_delay_6_mul_9_56
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_56_opA.fifo),
        .read_port(rd_mul_9_56_opA.fifo)
        );

	//add_18_6<->delay_7
	fifo_ms #(18,DEPTH,FLUX) fifo_add_18_6_delay_7
	(
	.clk(clk),
	.rst(rst),
	.write_port(wr_add_18_6_sum.fifo),
	.read_port(rd_delay_7_in_pel.fifo)
	);

//blocco bordo arancione fifo nel ppt

	//delay_7<->remove_h
	fifo_ms #(18,DEPTH,FLUX) fifo_delay_7_remove_h_0
	(
	.clk(clk),
	.rst(rst),
	.write_port(wr_delay_7_out_pel.fifo),
	.read_port(rd_remove_h_0_in_pel.fifo)
	);
	
	//add_18_13<->remove_h
	fifo_ms #(18,DEPTH,FLUX) fifo_add_18_13_remove_h_1
	(
	.clk(clk),
	.rst(rst),
	.write_port(wr_add_18_13_sum.fifo),
	.read_port(rd_remove_h_1_in_pel.fifo)
	);

	//add_18_20<->remove_h
	fifo_ms #(18,DEPTH,FLUX) fifo_add_18_20_remove_h_2
	(
	.clk(clk),
	.rst(rst),
	.write_port(wr_add_18_20_sum.fifo),
	.read_port(rd_remove_h_2_in_pel.fifo)
	);

	//add_18_27<->remove_h
	fifo_ms #(18,DEPTH,FLUX) fifo_add_18_27_remove_h_3
	(
	.clk(clk),
	.rst(rst),
	.write_port(wr_add_18_27_sum.fifo),
	.read_port(rd_remove_h_3_in_pel.fifo)
	);

	//add_18_34<->remove_h
	fifo_ms #(18,DEPTH,FLUX) fifo_add_18_34_remove_h_4
	(
	.clk(clk),
	.rst(rst),
	.write_port(wr_add_18_34_sum.fifo),
	.read_port(rd_remove_h_4_in_pel.fifo)
	);
	
	//add_18_41<->remove_h
	fifo_ms #(18,DEPTH,FLUX) fifo_add_18_41_remove_h_5
	(
	.clk(clk),
	.rst(rst),
	.write_port(wr_add_18_41_sum.fifo),
	.read_port(rd_remove_h_5_in_pel.fifo)
	);

	//add_18_48<->remove_h
	fifo_ms #(18,DEPTH,FLUX) fifo_add_18_48_remove_h_6
	(
	.clk(clk),
	.rst(rst),
	.write_port(wr_add_18_48_sum.fifo),
	.read_port(rd_remove_h_6_in_pel.fifo)
	);

	//add_18_55<->remove_h
	fifo_ms #(18,DEPTH,FLUX) fifo_add_18_55_remove_h_7
	(
	.clk(clk),
	.rst(rst),
	.write_port(wr_add_18_55_sum.fifo),
	.read_port(rd_remove_h_7_in_pel.fifo)
	);

        
   //coeff_h<->mul9 
    
    //1�riga 

        //coeff_luma_h<->mul_9_0
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_0_opB.fifo),
        .read_port(rd_mul_9_0_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_1
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_1_opB.fifo),
        .read_port(rd_mul_9_1_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_2
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_2_opB.fifo),
        .read_port(rd_mul_9_2_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_3
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_3_opB.fifo),
        .read_port(rd_mul_9_3_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_4
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_4_opB.fifo),
        .read_port(rd_mul_9_4_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_5
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_5_opB.fifo),
        .read_port(rd_mul_9_5_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_6
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_6_opB.fifo),
        .read_port(rd_mul_9_6_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_7
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_7_opB.fifo),
        .read_port(rd_mul_9_7_opB.fifo)
        );    
    
    //2� riga
    
        //coeff_luma_h<->mul_9_8
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_8
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_8_opB.fifo),
        .read_port(rd_mul_9_8_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_9
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_9
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_9_opB.fifo),
        .read_port(rd_mul_9_9_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_10
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_10
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_10_opB.fifo),
        .read_port(rd_mul_9_10_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_11
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_11
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_11_opB.fifo),
        .read_port(rd_mul_9_11_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_12
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_12
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_12_opB.fifo),
        .read_port(rd_mul_9_12_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_13
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_13
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_13_opB.fifo),
        .read_port(rd_mul_9_13_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_14
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_14
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_14_opB.fifo),
        .read_port(rd_mul_9_14_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_15
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_15
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_15_opB.fifo),
        .read_port(rd_mul_9_15_opB.fifo)
        );        
    
    //3� riga
    
        //coeff_luma_h<->mul_9_16
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_16
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_16_opB.fifo),
        .read_port(rd_mul_9_16_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_17
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_17
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_17_opB.fifo),
        .read_port(rd_mul_9_17_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_18
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_18
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_18_opB.fifo),
        .read_port(rd_mul_9_18_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_19
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_19
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_19_opB.fifo),
        .read_port(rd_mul_9_19_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_20
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_20
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_20_opB.fifo),
        .read_port(rd_mul_9_20_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_21
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_21
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_21_opB.fifo),
        .read_port(rd_mul_9_21_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_22
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_22
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_22_opB.fifo),
        .read_port(rd_mul_9_22_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_23
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_23
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_23_opB.fifo),
        .read_port(rd_mul_9_23_opB.fifo)
        );
            
    //4� riga
    
        //coeff_luma_h<->mul_9_24
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_24
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_24_opB.fifo),
        .read_port(rd_mul_9_24_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_25
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_25
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_25_opB.fifo),
        .read_port(rd_mul_9_25_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_26
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_26
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_26_opB.fifo),
        .read_port(rd_mul_9_26_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_27
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_27
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_27_opB.fifo),
        .read_port(rd_mul_9_27_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_28
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_28
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_28_opB.fifo),
        .read_port(rd_mul_9_28_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_29
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_29
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_29_opB.fifo),
        .read_port(rd_mul_9_29_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_30
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_30
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_30_opB.fifo),
        .read_port(rd_mul_9_30_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_31
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_31
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_31_opB.fifo),
        .read_port(rd_mul_9_31_opB.fifo)
        );
    
    //5� riga
    
        //coeff_luma_h<->mul_9_32
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_32
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_32_opB.fifo),
        .read_port(rd_mul_9_32_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_33
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_33
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_33_opB.fifo),
        .read_port(rd_mul_9_33_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_34
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_34
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_34_opB.fifo),
        .read_port(rd_mul_9_34_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_35
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_35
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_35_opB.fifo),
        .read_port(rd_mul_9_35_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_36
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_36
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_36_opB.fifo),
        .read_port(rd_mul_9_36_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_37
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_37
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_37_opB.fifo),
        .read_port(rd_mul_9_37_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_38
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_38
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_38_opB.fifo),
        .read_port(rd_mul_9_38_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_39
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_39
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_39_opB.fifo),
        .read_port(rd_mul_9_39_opB.fifo)
        );
    
    //6� riga
    
        //coeff_luma_h<->mul_9_40
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_40
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_40_opB.fifo),
        .read_port(rd_mul_9_40_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_41
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_41
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_41_opB.fifo),
        .read_port(rd_mul_9_41_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_42
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_42
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_42_opB.fifo),
        .read_port(rd_mul_9_42_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_43
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_43
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_43_opB.fifo),
        .read_port(rd_mul_9_43_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_44
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_44
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_44_opB.fifo),
        .read_port(rd_mul_9_44_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_45
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_45
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_45_opB.fifo),
        .read_port(rd_mul_9_45_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_46
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_46
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_46_opB.fifo),
        .read_port(rd_mul_9_46_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_47
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_47
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_47_opB.fifo),
        .read_port(rd_mul_9_47_opB.fifo)
        );
        
    //7� riga
    
        //coeff_luma_h<->mul_9_48
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_48
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_48_opB.fifo),
        .read_port(rd_mul_9_48_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_49
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_49
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_49_opB.fifo),
        .read_port(rd_mul_9_49_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_50
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_50
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_50_opB.fifo),
        .read_port(rd_mul_9_50_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_51
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_51
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_51_opB.fifo),
        .read_port(rd_mul_9_51_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_52
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_52
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_52_opB.fifo),
        .read_port(rd_mul_9_52_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_53
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_53
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_53_opB.fifo),
        .read_port(rd_mul_9_53_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_54
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_54
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_54_opB.fifo),
        .read_port(rd_mul_9_54_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_55
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_55
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_55_opB.fifo),
        .read_port(rd_mul_9_55_opB.fifo)
        );
            
    //8�riga
        
        //coeff_luma_h<->mul_9_56
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_56
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_56_opB.fifo),
        .read_port(rd_mul_9_56_opB.fifo)
        );        
        
        //coeff_luma_h<->mul_9_57
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_57
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_57_opB.fifo),
        .read_port(rd_mul_9_57_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_58
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_58
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_58_opB.fifo),
        .read_port(rd_mul_9_58_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_59
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_59
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_59_opB.fifo),
        .read_port(rd_mul_9_59_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_60
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_60
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_60_opB.fifo),
        .read_port(rd_mul_9_60_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_61
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_61
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_61_opB.fifo),
        .read_port(rd_mul_9_61_opB.fifo)
        );
        
        //coeff_luma_h<->mul_9_62
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_62
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_62_opB.fifo),
        .read_port(rd_mul_9_62_opB.fifo)
        );        

        //coeff_luma_h<->mul_9_63
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_h_mul_9_63
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_9_63_opB.fifo),
        .read_port(rd_mul_9_63_opB.fifo)
        );        

    //blocco bordo rosso fifo nel ppt
        
    //1� adder tree
        //mul_9_0<->adder_18_0
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_0_add_18_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_0_prod.fifo),
        .read_port(rd_add_18_0_opA.fifo)
        );

        //mul_9_1<->adder_18_0
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_1_add_18_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_1_prod.fifo),
        .read_port(rd_add_18_0_opB.fifo)
        );
        
        //mul_9_2<->adder_18_1
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_2_add_18_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_2_prod.fifo),
        .read_port(rd_add_18_1_opA.fifo)
        );  

        //mul_9_3<->adder_18_1
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_3_add_18_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_3_prod.fifo),
        .read_port(rd_add_18_1_opB.fifo)
        );

        //mul_9_4<->adder_18_2
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_4_add_18_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_4_prod.fifo),
        .read_port(rd_add_18_2_opA.fifo)
        );
        
        //mul_9_5<->adder_18_2
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_5_add_18_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_5_prod.fifo),
        .read_port(rd_add_18_2_opB.fifo)
        );

        //mul_9_6<->adder_18_3
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_6_add_18_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_6_prod.fifo),
        .read_port(rd_add_18_3_opA.fifo)
        );
        
        //mul_9_7<->adder_18_3
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_7_add_18_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_7_prod.fifo),
        .read_port(rd_add_18_3_opB.fifo)
        );

        //adder_18_0<->adder_18_4
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_0_add_18_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_0_sum.fifo),
        .read_port(rd_add_18_4_opA.fifo)
        );  

        //adder_18_1<->adder_18_4
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_1_add_18_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_1_sum.fifo),
        .read_port(rd_add_18_4_opB.fifo)
        );

        //adder_18_2<->adder_18_5
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_2_add_18_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_2_sum.fifo),
        .read_port(rd_add_18_5_opA.fifo)
        );
        
        //adder_18_3<->adder_18_5
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_3_add_18_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_3_sum.fifo),
        .read_port(rd_add_18_5_opB.fifo)
        );

        //adder_18_4<->adder_18_6
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_4_add_18_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_4_sum.fifo),
        .read_port(rd_add_18_6_opA.fifo)
        );
        
        //adder_18_5<->adder_18_6
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_5_add_18_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_5_sum.fifo),
        .read_port(rd_add_18_6_opB.fifo)
        );

    
    //2� adder tree

        //mul_9_8<->adder_18_7
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_8_add_18_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_8_prod.fifo),
        .read_port(rd_add_18_7_opA.fifo)
        );

        //mul_9_9<->adder_18_7
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_9_add_18_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_9_prod.fifo),
        .read_port(rd_add_18_7_opB.fifo)
        );
        
        //mul_9_10<->adder_18_8
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_10_9_add_18_8
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_10_prod.fifo),
        .read_port(rd_add_18_8_opA.fifo)
        );  

        //mul_9_11<->adder_18_8
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_11_add_18_8
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_11_prod.fifo),
        .read_port(rd_add_18_8_opB.fifo)
        );

        //mul_9_12<->adder_18_9
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_12_add_18_9
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_12_prod.fifo),
        .read_port(rd_add_18_9_opA.fifo)
        );
        
        //mul_9_13<->adder_18_9
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_13_add_18_9
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_13_prod.fifo),
        .read_port(rd_add_18_9_opB.fifo)
        );

        //mul_9_14<->adder_18_10
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_14_add_18_10
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_14_prod.fifo),
        .read_port(rd_add_18_10_opA.fifo)
        );
        
        //mul_9_15<->adder_18_10
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_15_add_18_10
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_15_prod.fifo),
        .read_port(rd_add_18_10_opB.fifo)
        );

        //adder_18_7<->adder_18_11
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_7_add_18_11
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_7_sum.fifo),
        .read_port(rd_add_18_11_opA.fifo)
        );  

        //adder_18_8<->adder_18_11
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_8_add_18_11
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_8_sum.fifo),
        .read_port(rd_add_18_11_opB.fifo)
        );

        //adder_18_9<->adder_18_12
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_9_add_18_12
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_9_sum.fifo),
        .read_port(rd_add_18_12_opA.fifo)
        );
        
        //adder_18_10<->adder_18_12
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_10_add_18_12
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_10_sum.fifo),
        .read_port(rd_add_18_12_opB.fifo)
        );

        //adder_18_11<->adder_18_13
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_11_add_18_13
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_11_sum.fifo),
        .read_port(rd_add_18_13_opA.fifo)
        );
        
        //adder_18_12<->adder_18_13
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_12_add_18_13
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_12_sum.fifo),
        .read_port(rd_add_18_13_opB.fifo)
        );
    
    //3� adder tree

        //mul_9_16<->adder_18_14
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_16_add_18_14
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_16_prod.fifo),
        .read_port(rd_add_18_14_opA.fifo)
        );

        //mul_9_17<->adder_18_14
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_17_add_18_14
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_17_prod.fifo),
        .read_port(rd_add_18_14_opB.fifo)
        );
        
        //mul_9_18<->adder_18_15
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_18_add_18_15
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_18_prod.fifo),
        .read_port(rd_add_18_15_opA.fifo)
        );  

        //mul_9_19<->adder_18_15
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_19_add_18_15
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_19_prod.fifo),
        .read_port(rd_add_18_15_opB.fifo)
        );

        //mul_9_20<->adder_18_16
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_20_add_18_16
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_20_prod.fifo),
        .read_port(rd_add_18_16_opA.fifo)
        );
        
        //mul_9_21<->adder_18_16
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_21_add_18_16
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_21_prod.fifo),
        .read_port(rd_add_18_16_opB.fifo)
        );

        //mul_9_22<->adder_18_17
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_22_add_18_17
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_22_prod.fifo),
        .read_port(rd_add_18_17_opA.fifo)
        );
        
        //mul_9_23<->adder_18_17
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_23_add_18_17
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_23_prod.fifo),
        .read_port(rd_add_18_17_opB.fifo)
        );

        //adder_18_14<->adder_18_18
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_14_add_18_18
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_14_sum.fifo),
        .read_port(rd_add_18_18_opA.fifo)
        );  

        //adder_18_15<->adder_18_18
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_15_add_18_18
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_15_sum.fifo),
        .read_port(rd_add_18_18_opB.fifo)
        );

        //adder_18_16<->adder_18_19
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_16_add_18_19
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_16_sum.fifo),
        .read_port(rd_add_18_19_opA.fifo)
        );
        
        //adder_18_17<->adder_18_19
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_17_add_18_19
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_17_sum.fifo),
        .read_port(rd_add_18_19_opB.fifo)
        );

        //adder_18_18<->adder_18_20
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_18_add_18_20
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_18_sum.fifo),
        .read_port(rd_add_18_20_opA.fifo)
        );
        
        //adder_18_19<->adder_18_20
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_19_add_18_20
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_19_sum.fifo),
        .read_port(rd_add_18_20_opB.fifo)
        );

    
    //4� adder tree

        //mul_9_24<->adder_18_21
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_24_add_18_21
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_24_prod.fifo),
        .read_port(rd_add_18_21_opA.fifo)
        );

        //mul_9_25<->adder_18_21
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_25_add_18_21
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_25_prod.fifo),
        .read_port(rd_add_18_21_opB.fifo)
        );
        
        //mul_9_26<->adder_18_22
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_26_add_18_22
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_26_prod.fifo),
        .read_port(rd_add_18_22_opA.fifo)
        );  

        //mul_9_27<->adder_18_22
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_27_add_18_22
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_27_prod.fifo),
        .read_port(rd_add_18_22_opB.fifo)
        );

        //mul_9_28<->adder_18_23
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_28_add_18_23
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_28_prod.fifo),
        .read_port(rd_add_18_23_opA.fifo)
        );
        
        //mul_9_29<->adder_18_23
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_29_add_18_23
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_29_prod.fifo),
        .read_port(rd_add_18_23_opB.fifo)
        );

        //mul_9_30<->adder_18_24
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_30_add_18_24
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_30_prod.fifo),
        .read_port(rd_add_18_24_opA.fifo)
        );
        
        //mul_9_31<->adder_18_24
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_31_add_18_24
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_31_prod.fifo),
        .read_port(rd_add_18_24_opB.fifo)
        );

        //adder_18_21<->adder_18_25
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_21_add_18_25
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_21_sum.fifo),
        .read_port(rd_add_18_25_opA.fifo)
        );  

        //adder_18_22<->adder_18_25
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_22_add_18_25
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_22_sum.fifo),
        .read_port(rd_add_18_25_opB.fifo)
        );

        //adder_18_23<->adder_18_26
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_23_add_18_26
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_23_sum.fifo),
        .read_port(rd_add_18_26_opA.fifo)
        );
        
        //adder_18_24<->adder_18_26
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_24_add_18_26
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_24_sum.fifo),
        .read_port(rd_add_18_26_opB.fifo)
        );

        //adder_18_25<->adder_18_27
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_25_add_18_27
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_25_sum.fifo),
        .read_port(rd_add_18_27_opA.fifo)
        );
        
        //adder_18_26<->adder_18_27
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_26_add_18_27
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_26_sum.fifo),
        .read_port(rd_add_18_27_opB.fifo)
        );
    
    //5� adder tree

        //mul_9_32<->adder_18_28
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_32_add_18_28
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_32_prod.fifo),
        .read_port(rd_add_18_28_opA.fifo)
        );

        //mul_9_33<->adder_18_28
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_33_add_18_28
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_33_prod.fifo),
        .read_port(rd_add_18_28_opB.fifo)
        );
        
        //mul_9_34<->adder_18_29
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_34_add_18_29
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_34_prod.fifo),
        .read_port(rd_add_18_29_opA.fifo)
        );  

        //mul_9_35<->adder_18_29
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_35_add_18_29
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_35_prod.fifo),
        .read_port(rd_add_18_29_opB.fifo)
        );

        //mul_9_36<->adder_18_30
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_36_add_18_30
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_36_prod.fifo),
        .read_port(rd_add_18_30_opA.fifo)
        );
        
        //mul_9_37<->adder_18_30
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_37_add_18_30
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_37_prod.fifo),
        .read_port(rd_add_18_30_opB.fifo)
        );

        //mul_9_38<->adder_18_31
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_38_add_18_31
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_38_prod.fifo),
        .read_port(rd_add_18_31_opA.fifo)
        );
        
        //mul_9_39<->adder_18_31
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_39_add_18_31
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_39_prod.fifo),
        .read_port(rd_add_18_31_opB.fifo)
        );

        //adder_18_28<->adder_18_32
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_28_add_18_32
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_28_sum.fifo),
        .read_port(rd_add_18_32_opA.fifo)
        );  

        //adder_18_29<->adder_18_32
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_29_add_18_32
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_29_sum.fifo),
        .read_port(rd_add_18_32_opB.fifo)
        );

        //adder_18_30<->adder_18_33
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_30_add_18_33
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_30_sum.fifo),
        .read_port(rd_add_18_33_opA.fifo)
        );
        
        //adder_18_31<->adder_18_33
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_31_add_18_33
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_31_sum.fifo),
        .read_port(rd_add_18_33_opB.fifo)
        );

        //adder_18_32<->adder_18_34
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_32_add_18_34
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_32_sum.fifo),
        .read_port(rd_add_18_34_opA.fifo)
        );
        
        //adder_18_33<->adder_18_34
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_33_add_18_34
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_33_sum.fifo),
        .read_port(rd_add_18_34_opB.fifo)
        );
    
    //6� adder tree

        //mul_9_40<->adder_18_35
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_40_add_18_35
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_40_prod.fifo),
        .read_port(rd_add_18_35_opA.fifo)
        );

        //mul_9_41<->adder_18_35
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_41_add_18_35
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_41_prod.fifo),
        .read_port(rd_add_18_35_opB.fifo)
        );
        
        //mul_9_42<->adder_18_36
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_42_add_18_36
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_42_prod.fifo),
        .read_port(rd_add_18_36_opA.fifo)
        );  

        //mul_9_43<->adder_18_36
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_43_add_18_36
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_43_prod.fifo),
        .read_port(rd_add_18_36_opB.fifo)
        );

        //mul_9_44<->adder_18_37
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_44_add_18_37
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_44_prod.fifo),
        .read_port(rd_add_18_37_opA.fifo)
        );
        
        //mul_9_45<->adder_18_37
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_45_add_18_37
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_45_prod.fifo),
        .read_port(rd_add_18_37_opB.fifo)
        );

        //mul_9_46<->adder_18_38
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_46_add_18_38
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_46_prod.fifo),
        .read_port(rd_add_18_38_opA.fifo)
        );
        
        //mul_9_47<->adder_18_38
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_47_add_18_38
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_47_prod.fifo),
        .read_port(rd_add_18_38_opB.fifo)
        );

        //adder_18_35<->adder_18_39
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_35_add_18_39
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_35_sum.fifo),
        .read_port(rd_add_18_39_opA.fifo)
        );  

        //adder_18_36<->adder_18_39
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_36_add_18_39
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_36_sum.fifo),
        .read_port(rd_add_18_39_opB.fifo)
        );

        //adder_18_37<->adder_18_40
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_37_add_18_40
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_37_sum.fifo),
        .read_port(rd_add_18_40_opA.fifo)
        );
        
        //adder_18_38<->adder_18_40
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_38_add_18_40
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_38_sum.fifo),
        .read_port(rd_add_18_40_opB.fifo)
        );

        //adder_18_39<->adder_18_41
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_39_add_18_41
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_39_sum.fifo),
        .read_port(rd_add_18_41_opA.fifo)
        );
        
        //adder_18_40<->adder_18_41
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_40_add_18_41
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_40_sum.fifo),
        .read_port(rd_add_18_41_opB.fifo)
        );
    
    //7� adder tree

        //mul_9_48<->adder_18_42
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_48_add_18_42
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_48_prod.fifo),
        .read_port(rd_add_18_42_opA.fifo)
        );

        //mul_9_49<->adder_18_42
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_49_add_18_42
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_49_prod.fifo),
        .read_port(rd_add_18_42_opB.fifo)
        );
        
        //mul_9_50<->adder_18_43
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_50_add_18_43
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_50_prod.fifo),
        .read_port(rd_add_18_43_opA.fifo)
        );  

        //mul_9_51<->adder_18_43
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_51_add_18_43
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_51_prod.fifo),
        .read_port(rd_add_18_43_opB.fifo)
        );

        //mul_9_52<->adder_18_44
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_52_add_18_44
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_52_prod.fifo),
        .read_port(rd_add_18_44_opA.fifo)
        );
        
        //mul_9_53<->adder_18_44
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_53_add_18_44
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_53_prod.fifo),
        .read_port(rd_add_18_44_opB.fifo)
        );

        //mul_9_54<->adder_18_45
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_54_add_18_45
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_54_prod.fifo),
        .read_port(rd_add_18_45_opA.fifo)
        );
        
        //mul_9_55<->adder_18_45
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_55_add_18_45
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_55_prod.fifo),
        .read_port(rd_add_18_45_opB.fifo)
        );

        //adder_18_42<->adder_18_46
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_42_add_18_46
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_42_sum.fifo),
        .read_port(rd_add_18_46_opA.fifo)
        );  

        //adder_18_43<->adder_18_46
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_43_add_18_46
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_43_sum.fifo),
        .read_port(rd_add_18_46_opB.fifo)
        );

        //adder_18_44<->adder_18_47
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_44_add_18_47
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_44_sum.fifo),
        .read_port(rd_add_18_47_opA.fifo)
        );
        
        //adder_18_45<->adder_18_47
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_45_add_18_47
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_45_sum.fifo),
        .read_port(rd_add_18_47_opB.fifo)
        );

        //adder_18_46<->adder_18_48
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_46_add_18_48
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_46_sum.fifo),
        .read_port(rd_add_18_48_opA.fifo)
        );
        
        //adder_18_47<->adder_18_48
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_47_add_18_48
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_47_sum.fifo),
        .read_port(rd_add_18_48_opB.fifo)
        );
    
    //8� adder tree       

        //mul_9_56<->adder_18_49
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_56_add_18_49
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_56_prod.fifo),
        .read_port(rd_add_18_49_opA.fifo)
        );

        //mul_9_57<->adder_18_49
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_57_add_18_49
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_57_prod.fifo),
        .read_port(rd_add_18_49_opB.fifo)
        );
        
        //mul_9_58<->adder_18_50
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_58_add_18_50
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_58_prod.fifo),
        .read_port(rd_add_18_50_opA.fifo)
        );  

        //mul_9_59<->adder_18_50
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_59_add_18_50
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_59_prod.fifo),
        .read_port(rd_add_18_50_opB.fifo)
        );

        //mul_9_60<->adder_18_51
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_60_add_18_51
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_60_prod.fifo),
        .read_port(rd_add_18_51_opA.fifo)
        );
        
        //mul_9_61<->adder_18_51
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_61_add_18_51
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_61_prod.fifo),
        .read_port(rd_add_18_51_opB.fifo)
        );

        //mul_9_62<->adder_18_52
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_62_add_18_52
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_62_prod.fifo),
        .read_port(rd_add_18_52_opA.fifo)
        );
        
        //mul_9_63<->adder_18_52
        fifo_ms #(18,DEPTH,FLUX) fifo_mul_9_63_add_18_52
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_9_63_prod.fifo),
        .read_port(rd_add_18_52_opB.fifo)
        );

        //adder_18_49<->adder_18_53
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_49_add_18_53
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_49_sum.fifo),
        .read_port(rd_add_18_53_opA.fifo)
        );  

        //adder_18_50<->adder_18_53
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_50_add_18_53
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_50_sum.fifo),
        .read_port(rd_add_18_53_opB.fifo)
        );

        //adder_18_51<->adder_18_54
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_51_add_18_54
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_51_sum.fifo),
        .read_port(rd_add_18_54_opA.fifo)
        );
        
        //adder_18_52<->adder_18_54
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_52_add_18_54
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_52_sum.fifo),
        .read_port(rd_add_18_54_opB.fifo)
        );

        //adder_18_53<->adder_18_55
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_53_add_18_55
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_53_sum.fifo),
        .read_port(rd_add_18_55_opA.fifo)
        );
        
        //adder_18_54<->adder_18_55
        fifo_ms #(18,DEPTH,FLUX) fifo_add_18_54_add_18_55
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_18_54_sum.fifo),
        .read_port(rd_add_18_55_opB.fifo)
        );


              
//FINE FIFO PRIMA PARTE



                      
//MODULI PRIMA PARTE



    //DELAY (x7); I: ORANGE - O: ORANGE / DARK YELLOW
     
        //delay0
        delay #(FLUX) delay_0 
        (
        .clk(clk),
        .rst(rst),
        .read_port_in_pel(rd_delay_0_in_pel.actor),
        .write_port_out_pel(wr_delay_0_out_pel.actor)        
        );
         
        //delay1 
        delay #(FLUX) delay_1 
        (
        .clk(clk),
        .rst(rst),
        .read_port_in_pel(rd_delay_1_in_pel.actor),
        .write_port_out_pel(wr_delay_1_out_pel.actor)        
        );    
        
        //delay2
        delay #(FLUX) delay_2 
        (
        .clk(clk),
        .rst(rst),
        .read_port_in_pel(rd_delay_2_in_pel.actor),
        .write_port_out_pel(wr_delay_2_out_pel.actor)        
        );
         
        //delay3 
        delay #(FLUX) delay_3 
        (
        .clk(clk),
        .rst(rst),
        .read_port_in_pel(rd_delay_3_in_pel.actor),
        .write_port_out_pel(wr_delay_3_out_pel.actor)        
        );    
    
        //delay4
        delay #(FLUX) delay_4 
        (
        .clk(clk),
        .rst(rst),
        .read_port_in_pel(rd_delay_4_in_pel.actor),
        .write_port_out_pel(wr_delay_4_out_pel.actor)        
        );
         
        //delay5 
        delay #(FLUX) delay_5 
        (
        .clk(clk),
        .rst(rst),
        .read_port_in_pel(rd_delay_5_in_pel.actor),
        .write_port_out_pel(wr_delay_5_out_pel.actor)        
        );    
    
        //delay6 
        delay #(FLUX) delay_6 
        (
        .clk(clk),
        .rst(rst),
        .read_port_in_pel(rd_delay_6_in_pel.actor),
        .write_port_out_pel(wr_delay_6_out_pel.actor)        
        );
		
        //delay7
        delay_d7 #(FLUX) delay_7 
        (
        .clk(clk),
        .rst(rst),
        .read_port_in_pel(rd_delay_7_in_pel.actor),
        .write_port_out_pel(wr_delay_7_out_pel.actor)        
        );		
				
    
    //COEFF_LUMA_H (x1); I: BLACK - O: BEIGE
    
        //coeff_luma_h
        coeff_luma #(FLUX) coeff_luma_h 
        (
        .read_port_alpha(rd_coeff_luma_h_alpha.actor),
        .write_port_c0(wr_coeff_luma_h_c0.actor),
        .write_port_c1(wr_coeff_luma_h_c1.actor),
        .write_port_c2(wr_coeff_luma_h_c2.actor),
        .write_port_c3(wr_coeff_luma_h_c3.actor),
        .write_port_c4(wr_coeff_luma_h_c4.actor),
        .write_port_c5(wr_coeff_luma_h_c5.actor),
        .write_port_c6(wr_coeff_luma_h_c6.actor),
        .write_port_c7(wr_coeff_luma_h_c7.actor)                               
        );    
    
        //COEFF_LUMA_V (x1); I: BLACK - O: GREEN (2�HALF)
        
        //coeff_luma_v
        coeff_luma #(FLUX) coeff_luma_v 
        (
        .read_port_alpha(rd_coeff_luma_v_alpha.actor),
        .write_port_c0(wr_coeff_luma_v_c0.actor),
        .write_port_c1(wr_coeff_luma_v_c1.actor),
        .write_port_c2(wr_coeff_luma_v_c2.actor),
        .write_port_c3(wr_coeff_luma_v_c3.actor),
        .write_port_c4(wr_coeff_luma_v_c4.actor),
        .write_port_c5(wr_coeff_luma_v_c5.actor),
        .write_port_c6(wr_coeff_luma_v_c6.actor),
        .write_port_c7(wr_coeff_luma_v_c7.actor)                               
        );

    //ADD18 (x56); I: BORDEAUX/GREEN - O: GREEN / YELLOW

	//1� adder tree
    
        //add18_0
        add_18 #(FLUX) add18_0
        (
        .read_port_opA(rd_add_18_0_opA.actor),
        .read_port_opB(rd_add_18_0_opB.actor),    
        .write_port_sum(wr_add_18_0_sum.actor)        
        );
    
        //add18_1 
        add_18 #(FLUX) add18_1 
        (
        .read_port_opA(rd_add_18_1_opA.actor),
        .read_port_opB(rd_add_18_1_opB.actor),    
        .write_port_sum(wr_add_18_1_sum.actor)        
        );
    
        //add18_2
        add_18 #(FLUX) add18_2 
        (
        .read_port_opA(rd_add_18_2_opA.actor),
        .read_port_opB(rd_add_18_2_opB.actor),    
        .write_port_sum(wr_add_18_2_sum.actor)        
        );
    
        //add18_3
        add_18 #(FLUX) add18_3
        (
        .read_port_opA(rd_add_18_3_opA.actor),
        .read_port_opB(rd_add_18_3_opB.actor),    
        .write_port_sum(wr_add_18_3_sum.actor)        
        );
        
        //add18_4 
        add_18 #(FLUX) add18_4 
        (
        .read_port_opA(rd_add_18_4_opA.actor),
        .read_port_opB(rd_add_18_4_opB.actor),    
        .write_port_sum(wr_add_18_4_sum.actor)        
        );
    
        //add18_5 
        add_18 #(FLUX) add18_5 
        (
        .read_port_opA(rd_add_18_5_opA.actor),
        .read_port_opB(rd_add_18_5_opB.actor),    
        .write_port_sum(wr_add_18_5_sum.actor)        
        );
        
        //add18_6
        add_18 #(FLUX) add18_6
        (
        .read_port_opA(rd_add_18_6_opA.actor),
        .read_port_opB(rd_add_18_6_opB.actor),    
        .write_port_sum(wr_add_18_6_sum.actor)        
        );

	//2� adder tree
    
        //add18_7
        add_18 #(FLUX) add18_7
        (
        .read_port_opA(rd_add_18_7_opA.actor),
        .read_port_opB(rd_add_18_7_opB.actor),    
        .write_port_sum(wr_add_18_7_sum.actor)        
        );
    
        //add18_8 
        add_18 #(FLUX) add18_8 
        (
        .read_port_opA(rd_add_18_8_opA.actor),
        .read_port_opB(rd_add_18_8_opB.actor),    
        .write_port_sum(wr_add_18_8_sum.actor)        
        );
    
        //add18_9
        add_18 #(FLUX) add18_9 
        (
        .read_port_opA(rd_add_18_9_opA.actor),
        .read_port_opB(rd_add_18_9_opB.actor),    
        .write_port_sum(wr_add_18_9_sum.actor)        
        );
    
        //add18_10
        add_18 #(FLUX) add18_10
        (
        .read_port_opA(rd_add_18_10_opA.actor),
        .read_port_opB(rd_add_18_10_opB.actor),    
        .write_port_sum(wr_add_18_10_sum.actor)        
        );
        
        //add18_11 
        add_18 #(FLUX) add18_11 
        (
        .read_port_opA(rd_add_18_11_opA.actor),
        .read_port_opB(rd_add_18_11_opB.actor),    
        .write_port_sum(wr_add_18_11_sum.actor)        
        );
    
        //add18_12 
        add_18 #(FLUX) add18_12
        (
        .read_port_opA(rd_add_18_12_opA.actor),
        .read_port_opB(rd_add_18_12_opB.actor),    
        .write_port_sum(wr_add_18_12_sum.actor)        
        );
        
        //add18_13
        add_18 #(FLUX) add18_13
        (
        .read_port_opA(rd_add_18_13_opA.actor),
        .read_port_opB(rd_add_18_13_opB.actor),    
        .write_port_sum(wr_add_18_13_sum.actor)        
        );
		
	//3� adder tree
    
        //add18_14
        add_18 #(FLUX) add18_14
        (
        .read_port_opA(rd_add_18_14_opA.actor),
        .read_port_opB(rd_add_18_14_opB.actor),    
        .write_port_sum(wr_add_18_14_sum.actor)        
        );
    
        //add18_15 
        add_18 #(FLUX) add18_15
        (
        .read_port_opA(rd_add_18_15_opA.actor),
        .read_port_opB(rd_add_18_15_opB.actor),    
        .write_port_sum(wr_add_18_15_sum.actor)        
        );
    
        //add18_16
        add_18 #(FLUX) add18_16
        (
        .read_port_opA(rd_add_18_16_opA.actor),
        .read_port_opB(rd_add_18_16_opB.actor),    
        .write_port_sum(wr_add_18_16_sum.actor)        
        );
    
        //add18_17
        add_18 #(FLUX) add18_17
        (
        .read_port_opA(rd_add_18_17_opA.actor),
        .read_port_opB(rd_add_18_17_opB.actor),    
        .write_port_sum(wr_add_18_17_sum.actor)        
        );
        
        //add18_18 
        add_18 #(FLUX) add18_18
        (
        .read_port_opA(rd_add_18_18_opA.actor),
        .read_port_opB(rd_add_18_18_opB.actor),    
        .write_port_sum(wr_add_18_18_sum.actor)        
        );
    
        //add18_19 
        add_18 #(FLUX) add18_19 
        (
        .read_port_opA(rd_add_18_19_opA.actor),
        .read_port_opB(rd_add_18_19_opB.actor),    
        .write_port_sum(wr_add_18_19_sum.actor)        
        );
        
        //add18_20
        add_18 #(FLUX) add18_20
        (
        .read_port_opA(rd_add_18_20_opA.actor),
        .read_port_opB(rd_add_18_20_opB.actor),    
        .write_port_sum(wr_add_18_20_sum.actor)        
        );		
		
	//4�adder tree
    
        //add18_21
        add_18 #(FLUX) add18_21
        (
        .read_port_opA(rd_add_18_21_opA.actor),
        .read_port_opB(rd_add_18_21_opB.actor),    
        .write_port_sum(wr_add_18_21_sum.actor)        
        );
    
        //add18_22
        add_18 #(FLUX) add18_22
        (
        .read_port_opA(rd_add_18_22_opA.actor),
        .read_port_opB(rd_add_18_22_opB.actor),    
        .write_port_sum(wr_add_18_22_sum.actor)        
        );
    
        //add18_23
        add_18 #(FLUX) add18_23
        (
        .read_port_opA(rd_add_18_23_opA.actor),
        .read_port_opB(rd_add_18_23_opB.actor),    
        .write_port_sum(wr_add_18_23_sum.actor)        
        );
    
        //add18_24
        add_18 #(FLUX) add18_24
        (
        .read_port_opA(rd_add_18_24_opA.actor),
        .read_port_opB(rd_add_18_24_opB.actor),    
        .write_port_sum(wr_add_18_24_sum.actor)        
        );
        
        //add18_25 
        add_18 #(FLUX) add18_25
        (
        .read_port_opA(rd_add_18_25_opA.actor),
        .read_port_opB(rd_add_18_25_opB.actor),    
        .write_port_sum(wr_add_18_25_sum.actor)        
        );
    
        //add18_26 
        add_18 #(FLUX) add18_26
        (
        .read_port_opA(rd_add_18_26_opA.actor),
        .read_port_opB(rd_add_18_26_opB.actor),    
        .write_port_sum(wr_add_18_26_sum.actor)        
        );
        
        //add18_27
        add_18 #(FLUX) add18_27
        (
        .read_port_opA(rd_add_18_27_opA.actor),
        .read_port_opB(rd_add_18_27_opB.actor),    
        .write_port_sum(wr_add_18_27_sum.actor)        
        );

	//5�adder tree
    
        //add18_28
        add_18 #(FLUX) add18_28
        (
        .read_port_opA(rd_add_18_28_opA.actor),
        .read_port_opB(rd_add_18_28_opB.actor),    
        .write_port_sum(wr_add_18_28_sum.actor)        
        );
    
        //add18_29
        add_18 #(FLUX) add18_29
        (
        .read_port_opA(rd_add_18_29_opA.actor),
        .read_port_opB(rd_add_18_29_opB.actor),    
        .write_port_sum(wr_add_18_29_sum.actor)        
        );
    
        //add18_30
        add_18 #(FLUX) add18_30
        (
        .read_port_opA(rd_add_18_30_opA.actor),
        .read_port_opB(rd_add_18_30_opB.actor),    
        .write_port_sum(wr_add_18_30_sum.actor)        
        );
    
        //add18_31
        add_18 #(FLUX) add18_31
        (
        .read_port_opA(rd_add_18_31_opA.actor),
        .read_port_opB(rd_add_18_31_opB.actor),    
        .write_port_sum(wr_add_18_31_sum.actor)        
        );
        
        //add18_32
        add_18 #(FLUX) add18_32
        (
        .read_port_opA(rd_add_18_32_opA.actor),
        .read_port_opB(rd_add_18_32_opB.actor),    
        .write_port_sum(wr_add_18_32_sum.actor)        
        );
    
        //add18_33
        add_18 #(FLUX) add18_33 
        (
        .read_port_opA(rd_add_18_33_opA.actor),
        .read_port_opB(rd_add_18_33_opB.actor),    
        .write_port_sum(wr_add_18_33_sum.actor)        
        );
        
        //add18_34
        add_18 #(FLUX) add18_34
        (
        .read_port_opA(rd_add_18_34_opA.actor),
        .read_port_opB(rd_add_18_34_opB.actor),    
        .write_port_sum(wr_add_18_34_sum.actor)        
        );

	//6�adder tree
    
        //add18_35
        add_18 #(FLUX) add18_35
        (
        .read_port_opA(rd_add_18_35_opA.actor),
        .read_port_opB(rd_add_18_35_opB.actor),    
        .write_port_sum(wr_add_18_35_sum.actor)        
        );
    
        //add18_36 
        add_18 #(FLUX) add18_36 
        (
        .read_port_opA(rd_add_18_36_opA.actor),
        .read_port_opB(rd_add_18_36_opB.actor),    
        .write_port_sum(wr_add_18_36_sum.actor)        
        );
    
        //add18_37
        add_18 #(FLUX) add18_37
        (
        .read_port_opA(rd_add_18_37_opA.actor),
        .read_port_opB(rd_add_18_37_opB.actor),    
        .write_port_sum(wr_add_18_37_sum.actor)        
        );
    
        //add18_38
        add_18 #(FLUX) add18_38
        (
        .read_port_opA(rd_add_18_38_opA.actor),
        .read_port_opB(rd_add_18_38_opB.actor),    
        .write_port_sum(wr_add_18_38_sum.actor)        
        );
        
        //add18_39 
        add_18 #(FLUX) add18_39
        (
        .read_port_opA(rd_add_18_39_opA.actor),
        .read_port_opB(rd_add_18_39_opB.actor),    
        .write_port_sum(wr_add_18_39_sum.actor)        
        );
    
        //add18_40 
        add_18 #(FLUX) add18_40
        (
        .read_port_opA(rd_add_18_40_opA.actor),
        .read_port_opB(rd_add_18_40_opB.actor),    
        .write_port_sum(wr_add_18_40_sum.actor)        
        );
        
        //add18_41
        add_18 #(FLUX) add18_41
        (
        .read_port_opA(rd_add_18_41_opA.actor),
        .read_port_opB(rd_add_18_41_opB.actor),    
        .write_port_sum(wr_add_18_41_sum.actor)        
        );
        
	//7�adder
    
        //add18_42
        add_18 #(FLUX) add18_42
        (
        .read_port_opA(rd_add_18_42_opA.actor),
        .read_port_opB(rd_add_18_42_opB.actor),    
        .write_port_sum(wr_add_18_42_sum.actor)        
        );
    
        //add18_43 
        add_18 #(FLUX) add18_43 
        (
        .read_port_opA(rd_add_18_43_opA.actor),
        .read_port_opB(rd_add_18_43_opB.actor),    
        .write_port_sum(wr_add_18_43_sum.actor)        
        );
    
        //add18_44
        add_18 #(FLUX) add18_44
        (
        .read_port_opA(rd_add_18_44_opA.actor),
        .read_port_opB(rd_add_18_44_opB.actor),    
        .write_port_sum(wr_add_18_44_sum.actor)        
        );
    
        //add18_45
        add_18 #(FLUX) add18_45
        (
        .read_port_opA(rd_add_18_45_opA.actor),
        .read_port_opB(rd_add_18_45_opB.actor),    
        .write_port_sum(wr_add_18_45_sum.actor)        
        );
        
        //add18_46 
        add_18 #(FLUX) add18_46 
        (
        .read_port_opA(rd_add_18_46_opA.actor),
        .read_port_opB(rd_add_18_46_opB.actor),    
        .write_port_sum(wr_add_18_46_sum.actor)        
        );
    
        //add18_47 
        add_18 #(FLUX) add18_47 
        (
        .read_port_opA(rd_add_18_47_opA.actor),
        .read_port_opB(rd_add_18_47_opB.actor),    
        .write_port_sum(wr_add_18_47_sum.actor)        
        );
        
        //add18_48
        add_18 #(FLUX) add18_48
        (
        .read_port_opA(rd_add_18_48_opA.actor),
        .read_port_opB(rd_add_18_48_opB.actor),    
        .write_port_sum(wr_add_18_48_sum.actor)        
        );

	//8� adder tree
    
        //add18_49
        add_18 #(FLUX) add18_49
        (
        .read_port_opA(rd_add_18_49_opA.actor),
        .read_port_opB(rd_add_18_49_opB.actor),    
        .write_port_sum(wr_add_18_49_sum.actor)        
        );
    
        //add18_50
        add_18 #(FLUX) add18_50 
        (
        .read_port_opA(rd_add_18_50_opA.actor),
        .read_port_opB(rd_add_18_50_opB.actor),    
        .write_port_sum(wr_add_18_50_sum.actor)        
        );
    
        //add18_51
        add_18 #(FLUX) add18_51
        (
        .read_port_opA(rd_add_18_51_opA.actor),
        .read_port_opB(rd_add_18_51_opB.actor),    
        .write_port_sum(wr_add_18_51_sum.actor)        
        );
    
        //add18_52
        add_18 #(FLUX) add18_52
        (
        .read_port_opA(rd_add_18_52_opA.actor),
        .read_port_opB(rd_add_18_52_opB.actor),    
        .write_port_sum(wr_add_18_52_sum.actor)        
        );
        
        //add18_53 
        add_18 #(FLUX) add18_53 
        (
        .read_port_opA(rd_add_18_53_opA.actor),
        .read_port_opB(rd_add_18_53_opB.actor),    
        .write_port_sum(wr_add_18_53_sum.actor)        
        );
    
        //add18_54 
        add_18 #(FLUX) add18_54 
        (
        .read_port_opA(rd_add_18_54_opA.actor),
        .read_port_opB(rd_add_18_54_opB.actor),    
        .write_port_sum(wr_add_18_54_sum.actor)        
        );
        
        //add18_55
        add_18 #(FLUX) add18_55
        (
        .read_port_opA(rd_add_18_55_opA.actor),
        .read_port_opB(rd_add_18_55_opB.actor),    
        .write_port_sum(wr_add_18_55_sum.actor)        
        );		
		
    //MUL9 (x64); I: DARK YELLOW/RED/BEIGE - O: BORDEAUX / GREEN
    
	//1� riga
	
        //mul9_0
        mul_9 #(FLUX) mul9_0
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_0_ext_size.actor),
        .read_port_opA(rd_mul_9_0_opA.actor),
        .read_port_opB(rd_mul_9_0_opB.actor),        
        .write_port_prod(wr_mul_9_0_prod.actor)        
        );
    
        //mul9_1
        mul_9 #(FLUX) mul9_1
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_1_ext_size.actor),
        .read_port_opA(rd_mul_9_1_opA.actor),
        .read_port_opB(rd_mul_9_1_opB.actor),        
        .write_port_prod(wr_mul_9_1_prod.actor)        
        );
    
        //mul9_2
        mul_9 #(FLUX) mul9_2
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_2_ext_size.actor),
        .read_port_opA(rd_mul_9_2_opA.actor),
        .read_port_opB(rd_mul_9_2_opB.actor),        
        .write_port_prod(wr_mul_9_2_prod.actor)        
        );
    
        //mul9_3
        mul_9 #(FLUX) mul9_3
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_3_ext_size.actor),
        .read_port_opA(rd_mul_9_3_opA.actor),
        .read_port_opB(rd_mul_9_3_opB.actor),        
        .write_port_prod(wr_mul_9_3_prod.actor)        
        );
    
        //mul9_4
        mul_9 #(FLUX) mul9_4
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_4_ext_size.actor),
        .read_port_opA(rd_mul_9_4_opA.actor),
        .read_port_opB(rd_mul_9_4_opB.actor),        
        .write_port_prod(wr_mul_9_4_prod.actor)        
        );
    
        //mul9_5
        mul_9 #(FLUX) mul9_5
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_5_ext_size.actor),
        .read_port_opA(rd_mul_9_5_opA.actor),
        .read_port_opB(rd_mul_9_5_opB.actor),        
        .write_port_prod(wr_mul_9_5_prod.actor)        
        );
    
        //mul9_6
        mul_9 #(FLUX) mul9_6
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_6_ext_size.actor),
        .read_port_opA(rd_mul_9_6_opA.actor),
        .read_port_opB(rd_mul_9_6_opB.actor),        
        .write_port_prod(wr_mul_9_6_prod.actor)        
        );
    
        //mul9_7
        mul_9 #(FLUX) mul9_7
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_7_ext_size.actor),
        .read_port_opA(rd_mul_9_7_opA.actor),
        .read_port_opB(rd_mul_9_7_opB.actor),        
        .write_port_prod(wr_mul_9_7_prod.actor)        
        );
    
	//2� riga

        //mul9_8
        mul_9 #(FLUX) mul9_8
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_8_ext_size.actor),
        .read_port_opA(rd_mul_9_8_opA.actor),
        .read_port_opB(rd_mul_9_8_opB.actor),        
        .write_port_prod(wr_mul_9_8_prod.actor)        
        );

        //mul9_9
        mul_9 #(FLUX) mul9_9
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_9_ext_size.actor),
        .read_port_opA(rd_mul_9_9_opA.actor),
        .read_port_opB(rd_mul_9_9_opB.actor),        
        .write_port_prod(wr_mul_9_9_prod.actor)        
        );
    
        //mul9_10
        mul_9 #(FLUX) mul9_10
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_10_ext_size.actor),
        .read_port_opA(rd_mul_9_10_opA.actor),
        .read_port_opB(rd_mul_9_10_opB.actor),        
        .write_port_prod(wr_mul_9_10_prod.actor)        
        );
    
        //mul9_11
        mul_9 #(FLUX) mul9_11
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_11_ext_size.actor),
        .read_port_opA(rd_mul_9_11_opA.actor),
        .read_port_opB(rd_mul_9_11_opB.actor),        
        .write_port_prod(wr_mul_9_11_prod.actor)        
        );
    
        //mul9_12
        mul_9 #(FLUX) mul9_12
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_12_ext_size.actor),
        .read_port_opA(rd_mul_9_12_opA.actor),
        .read_port_opB(rd_mul_9_12_opB.actor),        
        .write_port_prod(wr_mul_9_12_prod.actor)        
        );
    
        //mul9_13
        mul_9 #(FLUX) mul9_13
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_13_ext_size.actor),
        .read_port_opA(rd_mul_9_13_opA.actor),
        .read_port_opB(rd_mul_9_13_opB.actor),        
        .write_port_prod(wr_mul_9_13_prod.actor)        
        );
    
        //mul9_14
        mul_9 #(FLUX) mul9_14
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_14_ext_size.actor),
        .read_port_opA(rd_mul_9_14_opA.actor),
        .read_port_opB(rd_mul_9_14_opB.actor),        
        .write_port_prod(wr_mul_9_14_prod.actor)        
        );
        
        //mul9_15
        mul_9 #(FLUX) mul9_15
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_15_ext_size.actor),
        .read_port_opA(rd_mul_9_15_opA.actor),
        .read_port_opB(rd_mul_9_15_opB.actor),        
        .write_port_prod(wr_mul_9_15_prod.actor)        
        );
		
	//3�riga

        //mul9_16
        mul_9 #(FLUX) mul9_16
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_16_ext_size.actor),
        .read_port_opA(rd_mul_9_16_opA.actor),
        .read_port_opB(rd_mul_9_16_opB.actor),        
        .write_port_prod(wr_mul_9_16_prod.actor)        
        );
    
        //mul9_17
        mul_9 #(FLUX) mul9_17
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_17_ext_size.actor),
        .read_port_opA(rd_mul_9_17_opA.actor),
        .read_port_opB(rd_mul_9_17_opB.actor),        
        .write_port_prod(wr_mul_9_17_prod.actor)        
        );
    
        //mul9_18
        mul_9 #(FLUX) mul9_18
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_18_ext_size.actor),
        .read_port_opA(rd_mul_9_18_opA.actor),
        .read_port_opB(rd_mul_9_18_opB.actor),        
        .write_port_prod(wr_mul_9_18_prod.actor)        
        );
    
        //mul9_19
        mul_9 #(FLUX) mul9_19
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_19_ext_size.actor),
        .read_port_opA(rd_mul_9_19_opA.actor),
        .read_port_opB(rd_mul_9_19_opB.actor),        
        .write_port_prod(wr_mul_9_19_prod.actor)        
        );
    
        //mul9_20
        mul_9 #(FLUX) mul9_20
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_20_ext_size.actor),
        .read_port_opA(rd_mul_9_20_opA.actor),
        .read_port_opB(rd_mul_9_20_opB.actor),        
        .write_port_prod(wr_mul_9_20_prod.actor)        
        );
    
        //mul9_21
        mul_9 #(FLUX) mul9_21
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_21_ext_size.actor),
        .read_port_opA(rd_mul_9_21_opA.actor),
        .read_port_opB(rd_mul_9_21_opB.actor),        
        .write_port_prod(wr_mul_9_21_prod.actor)        
        );
    
        //mul9_22
        mul_9 #(FLUX) mul9_22
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_22_ext_size.actor),
        .read_port_opA(rd_mul_9_22_opA.actor),
        .read_port_opB(rd_mul_9_22_opB.actor),        
        .write_port_prod(wr_mul_9_22_prod.actor)        
        );
    
        //mul9_23
        mul_9 #(FLUX) mul9_23
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_23_ext_size.actor),
        .read_port_opA(rd_mul_9_23_opA.actor),
        .read_port_opB(rd_mul_9_23_opB.actor),        
        .write_port_prod(wr_mul_9_23_prod.actor)        
        );
		
	//4�riga

        //mul9_24
        mul_9 #(FLUX) mul9_24
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_24_ext_size.actor),
        .read_port_opA(rd_mul_9_24_opA.actor),
        .read_port_opB(rd_mul_9_24_opB.actor),        
        .write_port_prod(wr_mul_9_24_prod.actor)        
        );
    
        //mul9_25
        mul_9 #(FLUX) mul9_25
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_25_ext_size.actor),
        .read_port_opA(rd_mul_9_25_opA.actor),
        .read_port_opB(rd_mul_9_25_opB.actor),        
        .write_port_prod(wr_mul_9_25_prod.actor)        
        );
    
        //mul9_26
        mul_9 #(FLUX) mul9_26
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_26_ext_size.actor),
        .read_port_opA(rd_mul_9_26_opA.actor),
        .read_port_opB(rd_mul_9_26_opB.actor),        
        .write_port_prod(wr_mul_9_26_prod.actor)        
        );
    
        //mul9_27
        mul_9 #(FLUX) mul9_27
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_27_ext_size.actor),
        .read_port_opA(rd_mul_9_27_opA.actor),
        .read_port_opB(rd_mul_9_27_opB.actor),        
        .write_port_prod(wr_mul_9_27_prod.actor)        
        );
    
        //mul9_28
        mul_9 #(FLUX) mul9_28
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_28_ext_size.actor),
        .read_port_opA(rd_mul_9_28_opA.actor),
        .read_port_opB(rd_mul_9_28_opB.actor),        
        .write_port_prod(wr_mul_9_28_prod.actor)        
        );
    
        //mul9_29
        mul_9 #(FLUX) mul9_29
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_29_ext_size.actor),
        .read_port_opA(rd_mul_9_29_opA.actor),
        .read_port_opB(rd_mul_9_29_opB.actor),        
        .write_port_prod(wr_mul_9_29_prod.actor)        
        );
    
        //mul9_30
        mul_9 #(FLUX) mul9_30
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_30_ext_size.actor),
        .read_port_opA(rd_mul_9_30_opA.actor),
        .read_port_opB(rd_mul_9_30_opB.actor),        
        .write_port_prod(wr_mul_9_30_prod.actor)        
        );
    
        //mul9_31
        mul_9 #(FLUX) mul9_31
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_31_ext_size.actor),
        .read_port_opA(rd_mul_9_31_opA.actor),
        .read_port_opB(rd_mul_9_31_opB.actor),        
        .write_port_prod(wr_mul_9_31_prod.actor)        
        );
		
	//5�riga

        //mul9_32
        mul_9 #(FLUX) mul9_32
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_32_ext_size.actor),
        .read_port_opA(rd_mul_9_32_opA.actor),
        .read_port_opB(rd_mul_9_32_opB.actor),        
        .write_port_prod(wr_mul_9_32_prod.actor)        
        );
    
        //mul9_33
        mul_9 #(FLUX) mul9_33
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_33_ext_size.actor),
        .read_port_opA(rd_mul_9_33_opA.actor),
        .read_port_opB(rd_mul_9_33_opB.actor),        
        .write_port_prod(wr_mul_9_33_prod.actor)        
        );
    
        //mul9_34
        mul_9 #(FLUX) mul9_34
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_34_ext_size.actor),
        .read_port_opA(rd_mul_9_34_opA.actor),
        .read_port_opB(rd_mul_9_34_opB.actor),        
        .write_port_prod(wr_mul_9_34_prod.actor)        
        );
    
        //mul9_35
        mul_9 #(FLUX) mul9_35
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_35_ext_size.actor),
        .read_port_opA(rd_mul_9_35_opA.actor),
        .read_port_opB(rd_mul_9_35_opB.actor),        
        .write_port_prod(wr_mul_9_35_prod.actor)        
        );
    
        //mul9_36
        mul_9 #(FLUX) mul9_36
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_36_ext_size.actor),
        .read_port_opA(rd_mul_9_36_opA.actor),
        .read_port_opB(rd_mul_9_36_opB.actor),        
        .write_port_prod(wr_mul_9_36_prod.actor)        
        );
    
        //mul9_37
        mul_9 #(FLUX) mul9_37
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_37_ext_size.actor),
        .read_port_opA(rd_mul_9_37_opA.actor),
        .read_port_opB(rd_mul_9_37_opB.actor),        
        .write_port_prod(wr_mul_9_37_prod.actor)        
        );
    
        //mul9_38
        mul_9 #(FLUX) mul9_38
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_38_ext_size.actor),
        .read_port_opA(rd_mul_9_38_opA.actor),
        .read_port_opB(rd_mul_9_38_opB.actor),        
        .write_port_prod(wr_mul_9_38_prod.actor)        
        );
    
        //mul9_39
        mul_9 #(FLUX) mul9_39
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_39_ext_size.actor),
        .read_port_opA(rd_mul_9_39_opA.actor),
        .read_port_opB(rd_mul_9_39_opB.actor),        
        .write_port_prod(wr_mul_9_39_prod.actor)        
        );
		
	//6�riga

        //mul9_40
        mul_9 #(FLUX) mul9_40
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_40_ext_size.actor),
        .read_port_opA(rd_mul_9_40_opA.actor),
        .read_port_opB(rd_mul_9_40_opB.actor),        
        .write_port_prod(wr_mul_9_40_prod.actor)        
        );
    
        //mul9_41
        mul_9 #(FLUX) mul9_41
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_41_ext_size.actor),
        .read_port_opA(rd_mul_9_41_opA.actor),
        .read_port_opB(rd_mul_9_41_opB.actor),        
        .write_port_prod(wr_mul_9_41_prod.actor)        
        );
    
        //mul9_42
        mul_9 #(FLUX) mul9_42
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_42_ext_size.actor),
        .read_port_opA(rd_mul_9_42_opA.actor),
        .read_port_opB(rd_mul_9_42_opB.actor),        
        .write_port_prod(wr_mul_9_42_prod.actor)        
        );
    
        //mul9_43
        mul_9 #(FLUX) mul9_43
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_43_ext_size.actor),
        .read_port_opA(rd_mul_9_43_opA.actor),
        .read_port_opB(rd_mul_9_43_opB.actor),        
        .write_port_prod(wr_mul_9_43_prod.actor)        
        );
    
        //mul9_44
        mul_9 #(FLUX) mul9_44
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_44_ext_size.actor),
        .read_port_opA(rd_mul_9_44_opA.actor),
        .read_port_opB(rd_mul_9_44_opB.actor),        
        .write_port_prod(wr_mul_9_44_prod.actor)        
        );
    
        //mul9_45
        mul_9 #(FLUX) mul9_45
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_45_ext_size.actor),
        .read_port_opA(rd_mul_9_45_opA.actor),
        .read_port_opB(rd_mul_9_45_opB.actor),        
        .write_port_prod(wr_mul_9_45_prod.actor)        
        );
    
        //mul9_46
        mul_9 #(FLUX) mul9_46
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_46_ext_size.actor),
        .read_port_opA(rd_mul_9_46_opA.actor),
        .read_port_opB(rd_mul_9_46_opB.actor),        
        .write_port_prod(wr_mul_9_46_prod.actor)        
        );
    
        //mul9_47
        mul_9 #(FLUX) mul9_47
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_47_ext_size.actor),
        .read_port_opA(rd_mul_9_47_opA.actor),
        .read_port_opB(rd_mul_9_47_opB.actor),        
        .write_port_prod(wr_mul_9_47_prod.actor)        
        );
		
	//7�riga

        //mul9_48
        mul_9 #(FLUX) mul9_48
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_48_ext_size.actor),
        .read_port_opA(rd_mul_9_48_opA.actor),
        .read_port_opB(rd_mul_9_48_opB.actor),        
        .write_port_prod(wr_mul_9_48_prod.actor)        
        );
    
        //mul9_49
        mul_9 #(FLUX) mul9_49
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_49_ext_size.actor),
        .read_port_opA(rd_mul_9_49_opA.actor),
        .read_port_opB(rd_mul_9_49_opB.actor),        
        .write_port_prod(wr_mul_9_49_prod.actor)        
        );
    
        //mul9_50
        mul_9 #(FLUX) mul9_50
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_50_ext_size.actor),
        .read_port_opA(rd_mul_9_50_opA.actor),
        .read_port_opB(rd_mul_9_50_opB.actor),        
        .write_port_prod(wr_mul_9_50_prod.actor)        
        );
    
        //mul9_51
        mul_9 #(FLUX) mul9_51
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_51_ext_size.actor),
        .read_port_opA(rd_mul_9_51_opA.actor),
        .read_port_opB(rd_mul_9_51_opB.actor),        
        .write_port_prod(wr_mul_9_51_prod.actor)        
        );
    
        //mul9_52
        mul_9 #(FLUX) mul9_52
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_52_ext_size.actor),
        .read_port_opA(rd_mul_9_52_opA.actor),
        .read_port_opB(rd_mul_9_52_opB.actor),        
        .write_port_prod(wr_mul_9_52_prod.actor)        
        );
    
        //mul9_53
        mul_9 #(FLUX) mul9_53
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_53_ext_size.actor),
        .read_port_opA(rd_mul_9_53_opA.actor),
        .read_port_opB(rd_mul_9_53_opB.actor),        
        .write_port_prod(wr_mul_9_53_prod.actor)        
        );
    
        //mul9_54
        mul_9 #(FLUX) mul9_54
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_54_ext_size.actor),
        .read_port_opA(rd_mul_9_54_opA.actor),
        .read_port_opB(rd_mul_9_54_opB.actor),        
        .write_port_prod(wr_mul_9_54_prod.actor)        
        );
    
        //mul9_55
        mul_9 #(FLUX) mul9_55
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_55_ext_size.actor),
        .read_port_opA(rd_mul_9_55_opA.actor),
        .read_port_opB(rd_mul_9_55_opB.actor),        
        .write_port_prod(wr_mul_9_55_prod.actor)        
        );
		
	//8�riga

        //mul9_56
        mul_9 #(FLUX) mul9_56
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_56_ext_size.actor),
        .read_port_opA(rd_mul_9_56_opA.actor),
        .read_port_opB(rd_mul_9_56_opB.actor),        
        .write_port_prod(wr_mul_9_56_prod.actor)        
        );
    
        //mul9_57
        mul_9 #(FLUX) mul9_57
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_57_ext_size.actor),
        .read_port_opA(rd_mul_9_57_opA.actor),
        .read_port_opB(rd_mul_9_57_opB.actor),        
        .write_port_prod(wr_mul_9_57_prod.actor)        
        );
    
        //mul9_58
        mul_9 #(FLUX) mul9_58
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_58_ext_size.actor),
        .read_port_opA(rd_mul_9_58_opA.actor),
        .read_port_opB(rd_mul_9_58_opB.actor),        
        .write_port_prod(wr_mul_9_58_prod.actor)        
        );
    
        //mul9_59
        mul_9 #(FLUX) mul9_59
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_59_ext_size.actor),
        .read_port_opA(rd_mul_9_59_opA.actor),
        .read_port_opB(rd_mul_9_59_opB.actor),        
        .write_port_prod(wr_mul_9_59_prod.actor)        
        );
    
        //mul9_60
        mul_9 #(FLUX) mul9_60
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_60_ext_size.actor),
        .read_port_opA(rd_mul_9_60_opA.actor),
        .read_port_opB(rd_mul_9_60_opB.actor),        
        .write_port_prod(wr_mul_9_60_prod.actor)        
        );
    
        //mul9_61
        mul_9 #(FLUX) mul9_61
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_61_ext_size.actor),
        .read_port_opA(rd_mul_9_61_opA.actor),
        .read_port_opB(rd_mul_9_61_opB.actor),        
        .write_port_prod(wr_mul_9_61_prod.actor)        
        );
    
        //mul9_62
        mul_9 #(FLUX) mul9_62
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_62_ext_size.actor),
        .read_port_opA(rd_mul_9_62_opA.actor),
        .read_port_opB(rd_mul_9_62_opB.actor),        
        .write_port_prod(wr_mul_9_62_prod.actor)        
        );
    
        //mul9_63
        mul_9 #(FLUX) mul9_63
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_mul_9_63_ext_size.actor),
        .read_port_opA(rd_mul_9_63_opA.actor),
        .read_port_opB(rd_mul_9_63_opB.actor),        
        .write_port_prod(wr_mul_9_63_prod.actor)        
        );	
	
	
    //REMOVE_H (x8); I: LIME/YELLOW - O: DARK GREY (2�HALF) / RED (2�HALF)

        //remove_h_0
        remove_h #(FLUX) remove_h_0
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_remove_h_0_ext_size.actor),
        .read_port_in_pel(rd_remove_h_0_in_pel.actor),
		.write_port_out_pel(wr_remove_h_0_out_pel.actor)
        );
		
		//remove_h_1
        remove_h #(FLUX) remove_h_1
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_remove_h_1_ext_size.actor),
        .read_port_in_pel(rd_remove_h_1_in_pel.actor),
		.write_port_out_pel(wr_remove_h_1_out_pel.actor)
        );
		
		//remove_h_2
        remove_h #(FLUX) remove_h_2
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_remove_h_2_ext_size.actor),
        .read_port_in_pel(rd_remove_h_2_in_pel.actor),
		.write_port_out_pel(wr_remove_h_2_out_pel.actor)
        );
		
		//remove_h_3
        remove_h #(FLUX) remove_h_3
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_remove_h_3_ext_size.actor),
        .read_port_in_pel(rd_remove_h_3_in_pel.actor),
		.write_port_out_pel(wr_remove_h_3_out_pel.actor)
        );
		
		//remove_h_4
        remove_h #(FLUX) remove_h_4
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_remove_h_4_ext_size.actor),
        .read_port_in_pel(rd_remove_h_4_in_pel.actor),
		.write_port_out_pel(wr_remove_h_4_out_pel.actor)
        );
		
		//remove_h_5
        remove_h #(FLUX) remove_h_5
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_remove_h_5_ext_size.actor),
        .read_port_in_pel(rd_remove_h_5_in_pel.actor),
		.write_port_out_pel(wr_remove_h_5_out_pel.actor)
        );
		
		//remove_h_6
        remove_h #(FLUX) remove_h_6
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_remove_h_6_ext_size.actor),
        .read_port_in_pel(rd_remove_h_6_in_pel.actor),
		.write_port_out_pel(wr_remove_h_6_out_pel.actor)
        );
		
		//remove_h_7
        remove_h #(FLUX) remove_h_7
        (
        .clk(clk),
        .rst(rst),
        .read_port_ext_size(rd_remove_h_7_ext_size.actor),
        .read_port_in_pel(rd_remove_h_7_in_pel.actor),
		.write_port_out_pel(wr_remove_h_7_out_pel.actor)
        );
    
    //DERIVE (x1); I: LIGHT BLUE - O: LIME (2�HALF) / BROWN (2�HALF) / ORANGE (2�HALF)

        //derive_real_size
        derive_real_size #(FLUX) derive_real_size
        (
        .read_port_ext_size(rd_derive_real_size_ext_size.actor),       
        .write_port_real_size(wr_derive_real_size_real_size.actor)        
        );



//FINE MODULI PRIMA APRTE




//FIFO SECONDA PARTE



    //VIOLET: INPUT INPEL SHIFT (x8)
        
        //add_27_6<->shift_0
        fifo_ms #(27,DEPTH,FLUX) fifo_add27_6_shift_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_6_sum.fifo),
        .read_port(rd_shift_0_in_pel.fifo)
        );        

        //add_27_13<->shift_1
        fifo_ms #(27,DEPTH,FLUX) fifo_add27_13_shift_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_13_sum.fifo),
        .read_port(rd_shift_1_in_pel.fifo)
        );
		
        //add_27_20<->shift_2
        fifo_ms #(27,DEPTH,FLUX) fifo_add27_20_shift_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_20_sum.fifo),
        .read_port(rd_shift_2_in_pel.fifo)
        );

        //add_27_27<->shift_3
        fifo_ms #(27,DEPTH,FLUX) fifo_add27_27_shift_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_27_sum.fifo),
        .read_port(rd_shift_3_in_pel.fifo)
        );		

        //add_27_34<->shift_4
        fifo_ms #(27,DEPTH,FLUX) fifo_add27_34_shift_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_34_sum.fifo),
        .read_port(rd_shift_4_in_pel.fifo)
        );
		
        //add_27_41<->shift_5
        fifo_ms #(27,DEPTH,FLUX) fifo_add27_41_shift_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_41_sum.fifo),
        .read_port(rd_shift_5_in_pel.fifo)
        );		
		
        //add_27_48<->shift_6
        fifo_ms #(27,DEPTH,FLUX) fifo_add27_27_shift_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_48_sum.fifo),
        .read_port(rd_shift_6_in_pel.fifo)
        );		

        //add_27_55<->shift_7
        fifo_ms #(27,DEPTH,FLUX) fifo_add27_34_shift_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_55_sum.fifo),
        .read_port(rd_shift_7_in_pel.fifo)
        );
		
    
    //FUCSIA: INPUT INPEL CLIP (x8)    
    
        //shift_0<->clip_0
        fifo_ms #(16,DEPTH,FLUX) fifo_shift_0_clip_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_shift_0_out_pel.fifo),
        .read_port(rd_clip_0_in_pel.fifo)
        );

        //shift_1<->clip_1
        fifo_ms #(16,DEPTH,FLUX) fifo_shift_1_clip_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_shift_1_out_pel.fifo),
        .read_port(rd_clip_1_in_pel.fifo)
        );

        //shift_2<->clip_2
        fifo_ms #(16,DEPTH,FLUX) fifo_shift_2_clip_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_shift_2_out_pel.fifo),
        .read_port(rd_clip_2_in_pel.fifo)
        );

        //shift_3<->clip_3
        fifo_ms #(16,DEPTH,FLUX) fifo_shift_3_clip_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_shift_3_out_pel.fifo),
        .read_port(rd_clip_3_in_pel.fifo)
        );

        //shift_4<->clip_4
        fifo_ms #(16,DEPTH,FLUX) fifo_shift_4_clip_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_shift_4_out_pel.fifo),
        .read_port(rd_clip_4_in_pel.fifo)
        );

        //shift_5<->clip_5
        fifo_ms #(16,DEPTH,FLUX) fifo_shift_5_clip_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_shift_5_out_pel.fifo),
        .read_port(rd_clip_5_in_pel.fifo)
        );

        //shift_6<->clip_6
        fifo_ms #(16,DEPTH,FLUX) fifo_shift_6_clip_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_shift_6_out_pel.fifo),
        .read_port(rd_clip_6_in_pel.fifo)
        );

        //shift_7<->clip_7
        fifo_ms #(16,DEPTH,FLUX) fifo_shift_7_clip_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_shift_7_out_pel.fifo),
        .read_port(rd_clip_7_in_pel.fifo)
        );    
	
    //BROWN: INPUT REALSIZE REMOVE V
    
        //derive_real_size<->remove_v_0
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_remove_v_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_0_real_size.fifo),
        .read_port(rd_remove_v_0_real_size.fifo)
        );
    
        //derive_real_size<->remove_v_1
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_remove_v_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_1_real_size.fifo),
        .read_port(rd_remove_v_1_real_size.fifo)
        );
    
        //derive_real_size<->remove_v_2
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_remove_v_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_2_real_size.fifo),
        .read_port(rd_remove_v_2_real_size.fifo)
        );
    
        //derive_real_size<->remove_v_3
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_remove_v_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_3_real_size.fifo),
        .read_port(rd_remove_v_3_real_size.fifo)
        );
    
        //derive_real_size<->remove_v_4
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_remove_v_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_4_real_size.fifo),
        .read_port(rd_remove_v_4_real_size.fifo)
        );

        //derive_real_size<->remove_v_5
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_remove_v_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_5_real_size.fifo),
        .read_port(rd_remove_v_5_real_size.fifo)
        );
    
        //derive_real_size<->remove_v_6
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_remove_v_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_6_real_size.fifo),
        .read_port(rd_remove_v_6_real_size.fifo)
        );

        //derive_real_size<->remove_v_7
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_remove_v_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_7_real_size.fifo),
        .read_port(rd_remove_v_7_real_size.fifo)
        );

	
    //BLUE: INPUT EXTSIZE REMOVE V
    
        //extsize<->remove_v_0
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_v_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_0_ext_size.fifo),
        .read_port(rd_remove_v_0_ext_size.fifo)
        );       

        //extsize<->remove_v_1
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_v_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_1_ext_size.fifo),
        .read_port(rd_remove_v_1_ext_size.fifo)
        );       

        //extsize<->remove_v_2
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_v_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_2_ext_size.fifo),
        .read_port(rd_remove_v_2_ext_size.fifo)
        );       

        //extsize<->remove_v_3
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_v_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_3_ext_size.fifo),
        .read_port(rd_remove_v_3_ext_size.fifo)
        );       

        //extsize<->remove_v_4
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_v_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_4_ext_size.fifo),
        .read_port(rd_remove_v_4_ext_size.fifo)
        );       

        //extsize<->remove_v_5
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_v_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_5_ext_size.fifo),
        .read_port(rd_remove_v_5_ext_size.fifo)
        );       

        //extsize<->remove_v_6
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_v_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_6_ext_size.fifo),
        .read_port(rd_remove_v_6_ext_size.fifo)
        );       

        //extsize<->remove_v_7
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_remove_v_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_remove_v_7_ext_size.fifo),
        .read_port(rd_remove_v_7_ext_size.fifo)
        );       
        
    //PINK: INPUT INPEL REMOVE V (x8)

        //clip_0<->remove_v
        fifo_ms #(8,DEPTH,FLUX) fifo_clip_0_remove_v
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_clip_0_out_pel.fifo),
        .read_port(rd_remove_v_0_in_pel.fifo)
        );
		
        //clip_1<->remove_v
        fifo_ms #(8,DEPTH,FLUX) fifo_clip_1_remove_v
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_clip_1_out_pel.fifo),
        .read_port(rd_remove_v_1_in_pel.fifo)
        );

        //clip_2<->remove_v
        fifo_ms #(8,DEPTH,FLUX) fifo_clip_2_remove_v
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_clip_2_out_pel.fifo),
        .read_port(rd_remove_v_2_in_pel.fifo)
        );
		
        //clip_3<->remove_v
        fifo_ms #(8,DEPTH,FLUX) fifo_clip_3_remove_v
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_clip_3_out_pel.fifo),
        .read_port(rd_remove_v_3_in_pel.fifo)
        );

        //clip_4<->remove_v
        fifo_ms #(8,DEPTH,FLUX) fifo_clip_4_remove_v
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_clip_4_out_pel.fifo),
        .read_port(rd_remove_v_4_in_pel.fifo)
        );
		
        //clip_5<->remove_v
        fifo_ms #(8,DEPTH,FLUX) fifo_clip_5_remove_v
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_clip_5_out_pel.fifo),
        .read_port(rd_remove_v_5_in_pel.fifo)
        );

        //clip_6<->remove_v
        fifo_ms #(8,DEPTH,FLUX) fifo_clip_6_remove_v
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_clip_6_out_pel.fifo),
        .read_port(rd_remove_v_6_in_pel.fifo)
        );
		
        //clip_7<->remove_v
        fifo_ms #(8,DEPTH,FLUX) fifo_clip_7_remove_v
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_clip_7_out_pel.fifo),
        .read_port(rd_remove_v_7_in_pel.fifo)
        );

    //extsize mul18

    //1� riga                 
        //extsize<->mul_18_0        
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_0_ext_size.fifo),
        .read_port(rd_mul_18_0_ext_size.fifo)
        );        
                
        //extsize<->mul_18_1
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_1_ext_size.fifo),
        .read_port(rd_mul_18_1_ext_size.fifo)
        );
                
        //extsize<->mul_18_2
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_2_ext_size.fifo),
        .read_port(rd_mul_18_2_ext_size.fifo)
        );
        
        //extsize<->mul_18_3
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_3_ext_size.fifo),
        .read_port(rd_mul_18_3_ext_size.fifo)
        );
                
        //extsize<->mul_18_4
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_4_ext_size.fifo),
        .read_port(rd_mul_18_4_ext_size.fifo)
        );
        
        //extsize<->mul_18_5
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_5_ext_size.fifo),
        .read_port(rd_mul_18_5_ext_size.fifo)
        );        
        
        //extsize<->mul_18_6
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_6_ext_size.fifo),
        .read_port(rd_mul_18_6_ext_size.fifo)
        );
                
        //extsize<->mul_18_7
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_7_ext_size.fifo),
        .read_port(rd_mul_18_7_ext_size.fifo)
        );
  
    //2�riga
                   
        //extsize<->mul_18_8        
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_8
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_8_ext_size.fifo),
        .read_port(rd_mul_18_8_ext_size.fifo)
        );        
                
        //extsize<->mul_18_9
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_9
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_9_ext_size.fifo),
        .read_port(rd_mul_18_9_ext_size.fifo)
        );
                
        //extsize<->mul_18_10
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_10
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_10_ext_size.fifo),
        .read_port(rd_mul_18_10_ext_size.fifo)
        );
        
        //extsize<->mul_18_11
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_11
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_11_ext_size.fifo),
        .read_port(rd_mul_18_11_ext_size.fifo)
        );
                
        //extsize<->mul_18_12
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_12
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_12_ext_size.fifo),
        .read_port(rd_mul_18_12_ext_size.fifo)
        );
        
        //extsize<->mul_18_13
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_13
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_13_ext_size.fifo),
        .read_port(rd_mul_18_13_ext_size.fifo)
        );        
        
        //extsize<->mul_18_14
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_14
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_14_ext_size.fifo),
        .read_port(rd_mul_18_14_ext_size.fifo)
        );
                
        //extsize<->mul_18_15
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_15
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_15_ext_size.fifo),
        .read_port(rd_mul_18_15_ext_size.fifo)
        );
  
    //3�riga
                 
        //extsize<->mul_18_16        
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_16
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_16_ext_size.fifo),
        .read_port(rd_mul_18_16_ext_size.fifo)
        );        
                
        //extsize<->mul_18_17
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_17
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_17_ext_size.fifo),
        .read_port(rd_mul_18_17_ext_size.fifo)
        );
                
        //extsize<->mul_18_18
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_18
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_18_ext_size.fifo),
        .read_port(rd_mul_18_18_ext_size.fifo)
        );
        
        //extsize<->mul_18_19
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_19
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_19_ext_size.fifo),
        .read_port(rd_mul_18_19_ext_size.fifo)
        );
                
        //extsize<->mul_18_20
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_20
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_20_ext_size.fifo),
        .read_port(rd_mul_18_20_ext_size.fifo)
        );
        
        //extsize<->mul_18_21
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_21
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_21_ext_size.fifo),
        .read_port(rd_mul_18_21_ext_size.fifo)
        );        
        
        //extsize<->mul_18_22
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_22
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_22_ext_size.fifo),
        .read_port(rd_mul_18_22_ext_size.fifo)
        );
                
        //extsize<->mul_18_23
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_23
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_23_ext_size.fifo),
        .read_port(rd_mul_18_23_ext_size.fifo)
        );
    
    //4�riga
                     
        //extsize<->mul_18_24        
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_24
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_24_ext_size.fifo),
        .read_port(rd_mul_18_24_ext_size.fifo)
        );        
                
        //extsize<->mul_18_25
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_25
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_25_ext_size.fifo),
        .read_port(rd_mul_18_25_ext_size.fifo)
        );
                
        //extsize<->mul_18_26
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_26
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_26_ext_size.fifo),
        .read_port(rd_mul_18_26_ext_size.fifo)
        );
        
        //extsize<->mul_18_27
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_27
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_27_ext_size.fifo),
        .read_port(rd_mul_18_27_ext_size.fifo)
        );
                
        //extsize<->mul_18_28
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_28
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_28_ext_size.fifo),
        .read_port(rd_mul_18_28_ext_size.fifo)
        );
        
        //extsize<->mul_18_29
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_29
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_29_ext_size.fifo),
        .read_port(rd_mul_18_29_ext_size.fifo)
        );        
        
        //extsize<->mul_18_30
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_30
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_30_ext_size.fifo),
        .read_port(rd_mul_18_30_ext_size.fifo)
        );
                
        //extsize<->mul_18_31
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_31
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_31_ext_size.fifo),
        .read_port(rd_mul_18_31_ext_size.fifo)
        );
            
    //5�riga

        //extsize<->mul_18_32
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_32
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_32_ext_size.fifo),
        .read_port(rd_mul_18_32_ext_size.fifo)
        );        
                
        //extsize<->mul_18_33
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_33
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_33_ext_size.fifo),
        .read_port(rd_mul_18_33_ext_size.fifo)
        );
                
        //extsize<->mul_18_34
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_34
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_34_ext_size.fifo),
        .read_port(rd_mul_18_34_ext_size.fifo)
        );
        
        //extsize<->mul_18_35
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_35
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_35_ext_size.fifo),
        .read_port(rd_mul_18_35_ext_size.fifo)
        );
                
        //extsize<->mul_18_36
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_36
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_36_ext_size.fifo),
        .read_port(rd_mul_18_36_ext_size.fifo)
        );
        
        //extsize<->mul_18_37
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_37
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_37_ext_size.fifo),
        .read_port(rd_mul_18_37_ext_size.fifo)
        );        
        
        //extsize<->mul_18_38
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_38
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_38_ext_size.fifo),
        .read_port(rd_mul_18_38_ext_size.fifo)
        );
                
        //extsize<->mul_18_39
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_39
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_39_ext_size.fifo),
        .read_port(rd_mul_18_39_ext_size.fifo)
        );
    
    //6�riga
        
        //extsize<->mul_18_40
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_40
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_40_ext_size.fifo),
        .read_port(rd_mul_18_40_ext_size.fifo)
        );        
                
        //extsize<->mul_18_41
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_41
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_41_ext_size.fifo),
        .read_port(rd_mul_18_41_ext_size.fifo)
        );
                
        //extsize<->mul_18_42
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_42
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_42_ext_size.fifo),
        .read_port(rd_mul_18_42_ext_size.fifo)
        );
        
        //extsize<->mul_18_43
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_43
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_43_ext_size.fifo),
        .read_port(rd_mul_18_43_ext_size.fifo)
        );
                
        //extsize<->mul_18_44
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_44
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_44_ext_size.fifo),
        .read_port(rd_mul_18_44_ext_size.fifo)
        );
        
        //extsize<->mul_18_45
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_45
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_45_ext_size.fifo),
        .read_port(rd_mul_18_45_ext_size.fifo)
        );        
        
        //extsize<->mul_18_46
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_46
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_46_ext_size.fifo),
        .read_port(rd_mul_18_46_ext_size.fifo)
        );
                
        //extsize<->mul_18_47
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_47
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_47_ext_size.fifo),
        .read_port(rd_mul_18_47_ext_size.fifo)
        );
    
    //7�riga
        
        //extsize<->mul_18_48
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_48
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_48_ext_size.fifo),
        .read_port(rd_mul_18_48_ext_size.fifo)
        );        
                
        //extsize<->mul_18_49
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_49
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_49_ext_size.fifo),
        .read_port(rd_mul_18_49_ext_size.fifo)
        );
                
        //extsize<->mul_18_50
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_50
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_50_ext_size.fifo),
        .read_port(rd_mul_18_50_ext_size.fifo)
        );
        
        //extsize<->mul_18_51
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_51
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_51_ext_size.fifo),
        .read_port(rd_mul_18_51_ext_size.fifo)
        );
                
        //extsize<->mul_18_52
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_52
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_52_ext_size.fifo),
        .read_port(rd_mul_18_52_ext_size.fifo)
        );
        
        //extsize<->mul_18_53
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_53
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_53_ext_size.fifo),
        .read_port(rd_mul_18_53_ext_size.fifo)
        );        
        
        //extsize<->mul_18_54
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_54
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_54_ext_size.fifo),
        .read_port(rd_mul_18_54_ext_size.fifo)
        );
                
        //extsize<->mul_18_55
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_55
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_55_ext_size.fifo),
        .read_port(rd_mul_18_55_ext_size.fifo)
        );    
    
    //8�riga
        
        //extsize<->mul_18_56
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_56
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_56_ext_size.fifo),
        .read_port(rd_mul_18_56_ext_size.fifo)
        );        
                
        //extsize<->mul_18_57
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_57
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_57_ext_size.fifo),
        .read_port(rd_mul_18_57_ext_size.fifo)
        );
                
        //extsize<->mul_18_58
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_58
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_58_ext_size.fifo),
        .read_port(rd_mul_18_58_ext_size.fifo)
        );
        
        //extsize<->mul_18_59
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_59
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_59_ext_size.fifo),
        .read_port(rd_mul_18_59_ext_size.fifo)
        );
                
        //extsize<->mul_18_60
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_60
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_60_ext_size.fifo),
        .read_port(rd_mul_18_60_ext_size.fifo)
        );
        
        //extsize<->mul_18_61
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_61
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_61_ext_size.fifo),
        .read_port(rd_mul_18_61_ext_size.fifo)
        );        
        
        //extsize<->mul_18_62
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_62
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_62_ext_size.fifo),
        .read_port(rd_mul_18_62_ext_size.fifo)
        );
                
        //extsize<->mul_18_63
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_mul18_63
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_63_ext_size.fifo),
        .read_port(rd_mul_18_63_ext_size.fifo)
        );
	
    //realsize mul18

    //1� riga                 
        //realsize<->mul_18_0        
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_0_real_size.fifo),
        .read_port(rd_mul_18_0_real_size.fifo)
        );        
                
        //realsize<->mul_18_1
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_1_real_size.fifo),
        .read_port(rd_mul_18_1_real_size.fifo)
        );
                
        //realsize<->mul_18_2
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_2_real_size.fifo),
        .read_port(rd_mul_18_2_real_size.fifo)
        );
        
        //realsize<->mul_18_3
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_3_real_size.fifo),
        .read_port(rd_mul_18_3_real_size.fifo)
        );
                
        //realsize<->mul_18_4
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_4_real_size.fifo),
        .read_port(rd_mul_18_4_real_size.fifo)
        );
        
        //realsize<->mul_18_5
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_5_real_size.fifo),
        .read_port(rd_mul_18_5_real_size.fifo)
        );        
        
        //realsize<->mul_18_6
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_6_real_size.fifo),
        .read_port(rd_mul_18_6_real_size.fifo)
        );
                
        //realsize<->mul_18_7
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_7_real_size.fifo),
        .read_port(rd_mul_18_7_real_size.fifo)
        );
  
    //2�riga
                   
        //realsize<->mul_18_8        
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_8
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_8_real_size.fifo),
        .read_port(rd_mul_18_8_real_size.fifo)
        );        
                
        //realsize<->mul_18_9
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_9
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_9_real_size.fifo),
        .read_port(rd_mul_18_9_real_size.fifo)
        );
                
        //realsize<->mul_18_10
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_10
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_10_real_size.fifo),
        .read_port(rd_mul_18_10_real_size.fifo)
        );
        
        //realsize<->mul_18_11
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_11
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_11_real_size.fifo),
        .read_port(rd_mul_18_11_real_size.fifo)
        );
                
        //realsize<->mul_18_12
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_12
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_12_real_size.fifo),
        .read_port(rd_mul_18_12_real_size.fifo)
        );
        
        //realsize<->mul_18_13
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_13
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_13_real_size.fifo),
        .read_port(rd_mul_18_13_real_size.fifo)
        );        
        
        //realsize<->mul_18_14
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_14
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_14_real_size.fifo),
        .read_port(rd_mul_18_14_real_size.fifo)
        );
                
        //realsize<->mul_18_15
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_15
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_15_real_size.fifo),
        .read_port(rd_mul_18_15_real_size.fifo)
        );
  
    //3�riga
                 
        //realsize<->mul_18_16        
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_16
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_16_real_size.fifo),
        .read_port(rd_mul_18_16_real_size.fifo)
        );        
                
        //realsize<->mul_18_17
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_17
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_17_real_size.fifo),
        .read_port(rd_mul_18_17_real_size.fifo)
        );
                
        //realsize<->mul_18_18
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_18
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_18_real_size.fifo),
        .read_port(rd_mul_18_18_real_size.fifo)
        );
        
        //realsize<->mul_18_19
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_19
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_19_real_size.fifo),
        .read_port(rd_mul_18_19_real_size.fifo)
        );
                
        //realsize<->mul_18_20
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_20
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_20_real_size.fifo),
        .read_port(rd_mul_18_20_real_size.fifo)
        );
        
        //realsize<->mul_18_21
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_21
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_21_real_size.fifo),
        .read_port(rd_mul_18_21_real_size.fifo)
        );        
        
        //realsize<->mul_18_22
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_22
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_22_real_size.fifo),
        .read_port(rd_mul_18_22_real_size.fifo)
        );
                
        //realsize<->mul_18_23
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_23
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_23_real_size.fifo),
        .read_port(rd_mul_18_23_real_size.fifo)
        );
    
    //4�riga
                     
        //realsize<->mul_18_24        
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_24
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_24_real_size.fifo),
        .read_port(rd_mul_18_24_real_size.fifo)
        );        
                
        //realsize<->mul_18_25
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_25
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_25_real_size.fifo),
        .read_port(rd_mul_18_25_real_size.fifo)
        );
                
        //realsize<->mul_18_26
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_26
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_26_real_size.fifo),
        .read_port(rd_mul_18_26_real_size.fifo)
        );
        
        //realsize<->mul_18_27
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_27
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_27_real_size.fifo),
        .read_port(rd_mul_18_27_real_size.fifo)
        );
                
        //realsize<->mul_18_28
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_28
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_28_real_size.fifo),
        .read_port(rd_mul_18_28_real_size.fifo)
        );
        
        //realsize<->mul_18_29
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_29
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_29_real_size.fifo),
        .read_port(rd_mul_18_29_real_size.fifo)
        );        
        
        //realsize<->mul_18_30
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_30
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_30_real_size.fifo),
        .read_port(rd_mul_18_30_real_size.fifo)
        );
                
        //realsize<->mul_18_31
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_31
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_31_real_size.fifo),
        .read_port(rd_mul_18_31_real_size.fifo)
        );
            
    //5�riga

        //realsize<->mul_18_32
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_32
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_32_real_size.fifo),
        .read_port(rd_mul_18_32_real_size.fifo)
        );        
                
        //realsize<->mul_18_33
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_33
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_33_real_size.fifo),
        .read_port(rd_mul_18_33_real_size.fifo)
        );
                
        //realsize<->mul_18_34
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_34
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_34_real_size.fifo),
        .read_port(rd_mul_18_34_real_size.fifo)
        );
        
        //realsize<->mul_18_35
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_35
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_35_real_size.fifo),
        .read_port(rd_mul_18_35_real_size.fifo)
        );
                
        //realsize<->mul_18_36
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_36
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_36_real_size.fifo),
        .read_port(rd_mul_18_36_real_size.fifo)
        );
        
        //realsize<->mul_18_37
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_37
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_37_real_size.fifo),
        .read_port(rd_mul_18_37_real_size.fifo)
        );        
        
        //realsize<->mul_18_38
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_38
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_38_real_size.fifo),
        .read_port(rd_mul_18_38_real_size.fifo)
        );
                
        //realsize<->mul_18_39
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_39
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_39_real_size.fifo),
        .read_port(rd_mul_18_39_real_size.fifo)
        );
    
    //6�riga
        
        //realsize<->mul_18_40
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_40
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_40_real_size.fifo),
        .read_port(rd_mul_18_40_real_size.fifo)
        );        
                
        //realsize<->mul_18_41
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_41
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_41_real_size.fifo),
        .read_port(rd_mul_18_41_real_size.fifo)
        );
                
        //realsize<->mul_18_42
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_42
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_42_real_size.fifo),
        .read_port(rd_mul_18_42_real_size.fifo)
        );
        
        //realsize<->mul_18_43
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_43
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_43_real_size.fifo),
        .read_port(rd_mul_18_43_real_size.fifo)
        );
                
        //realsize<->mul_18_44
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_44
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_44_real_size.fifo),
        .read_port(rd_mul_18_44_real_size.fifo)
        );
        
        //realsize<->mul_18_45
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_45
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_45_real_size.fifo),
        .read_port(rd_mul_18_45_real_size.fifo)
        );        
        
        //realsize<->mul_18_46
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_46
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_46_real_size.fifo),
        .read_port(rd_mul_18_46_real_size.fifo)
        );
                
        //realsize<->mul_18_47
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_47
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_47_real_size.fifo),
        .read_port(rd_mul_18_47_real_size.fifo)
        );
    
    //7�riga
        
        //realsize<->mul_18_48
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_48
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_48_real_size.fifo),
        .read_port(rd_mul_18_48_real_size.fifo)
        );        
                
        //realsize<->mul_18_49
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_49
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_49_real_size.fifo),
        .read_port(rd_mul_18_49_real_size.fifo)
        );
                
        //realsize<->mul_18_50
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_50
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_50_real_size.fifo),
        .read_port(rd_mul_18_50_real_size.fifo)
        );
        
        //realsize<->mul_18_51
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_51
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_51_real_size.fifo),
        .read_port(rd_mul_18_51_real_size.fifo)
        );
                
        //realsize<->mul_18_52
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_52
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_52_real_size.fifo),
        .read_port(rd_mul_18_52_real_size.fifo)
        );
        
        //realsize<->mul_18_53
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_53
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_53_real_size.fifo),
        .read_port(rd_mul_18_53_real_size.fifo)
        );        
        
        //realsize<->mul_18_54
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_54
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_54_real_size.fifo),
        .read_port(rd_mul_18_54_real_size.fifo)
        );
                
        //realsize<->mul_18_55
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_55
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_55_real_size.fifo),
        .read_port(rd_mul_18_55_real_size.fifo)
        );    
    
    //8�riga
        
        //realsize<->mul_18_56
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_56
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_56_real_size.fifo),
        .read_port(rd_mul_18_56_real_size.fifo)
        );        
                
        //realsize<->mul_18_57
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_57
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_57_real_size.fifo),
        .read_port(rd_mul_18_57_real_size.fifo)
        );
                
        //realsize<->mul_18_58
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_58
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_58_real_size.fifo),
        .read_port(rd_mul_18_58_real_size.fifo)
        );
        
        //realsize<->mul_18_59
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_59
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_59_real_size.fifo),
        .read_port(rd_mul_18_59_real_size.fifo)
        );
                
        //realsize<->mul_18_60
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_60
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_60_real_size.fifo),
        .read_port(rd_mul_18_60_real_size.fifo)
        );
        
        //realsize<->mul_18_61
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_61
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_61_real_size.fifo),
        .read_port(rd_mul_18_61_real_size.fifo)
        );        
        
        //realsize<->mul_18_62
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_62
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_62_real_size.fifo),
        .read_port(rd_mul_18_62_real_size.fifo)
        );
                
        //realsize<->mul_18_63
        fifo_ms #(7,DEPTH,FLUX) fifo_realsize_mul18_63
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_63_real_size.fifo),
        .read_port(rd_mul_18_63_real_size.fifo)
        );	
	
	//Blocco celeste fifo nel ppt
   
	//1� colonna
   
        //remove_h0<->mul18_0
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_0_mul_18_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_0_opA.fifo),
        .read_port(rd_mul_18_0_opA.fifo)
        );

        //line_buffer0<->mul18_1
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_0_mul_18_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_1_opA.fifo),
        .read_port(rd_mul_18_1_opA.fifo)
        );

        //line_buffer_1<->mul18_2
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_0_mul_18_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_2_opA.fifo),
        .read_port(rd_mul_18_2_opA.fifo)
        );

        //line_buffer_2<->mul18_3
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_0_mul_18_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_3_opA.fifo),
        .read_port(rd_mul_18_3_opA.fifo)
        );

        //line_buffer_3<->mul18_4
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_0_mul_18_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_4_opA.fifo),
        .read_port(rd_mul_18_4_opA.fifo)
        );

        //line_buffer_4<->mul18_5
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_0_mul_18_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_5_opA.fifo),
        .read_port(rd_mul_18_5_opA.fifo)
        );

        //line_buffer_5<->mul18_6
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_0_mul_18_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_6_opA.fifo),
        .read_port(rd_mul_18_6_opA.fifo)
        );

        //line_buffer_6<->mul18_7
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_6_0_mul_18_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_line_buffer_6_0_out_pel.fifo),
        .read_port(rd_mul_18_7_opA.fifo)
        );

	//2� colonna
        
        //remove_h1<->mul18_8
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_1_mul_18_8
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_8_opA.fifo),
        .read_port(rd_mul_18_8_opA.fifo)
        );
                      
        //line_buffer_0<->mul18_9
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_1_mul_18_9
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_9_opA.fifo),
        .read_port(rd_mul_18_9_opA.fifo)
        );        
 
        //line_buffer_1<->mul18_10
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_1_mul_18_10
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_10_opA.fifo),
        .read_port(rd_mul_18_10_opA.fifo)
        );

        //line_buffer_2<->mul18_11
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_1_mul_18_11
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_11_opA.fifo),
        .read_port(rd_mul_18_11_opA.fifo)
        );        

        //line_buffer_3<->mul18_12
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_1_mul_18_12
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_12_opA.fifo),
        .read_port(rd_mul_18_12_opA.fifo)
        );        

        //line_buffer_4<->mul18_13
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_1_mul_18_13
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_13_opA.fifo),
        .read_port(rd_mul_18_13_opA.fifo)
        );      
 
         //line_buffer_5<->mul18_14
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_1_mul_18_14
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_14_opA.fifo),
        .read_port(rd_mul_18_14_opA.fifo)
        );      
 
         //line_buffer_6<->mul18_15
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_6_1_mul_18_15
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_line_buffer_6_1_out_pel.fifo),
        .read_port(rd_mul_18_15_opA.fifo)
        );      
 
	//3�colonna
    
        //remove_h2<->mul18_16
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_2_mul_18_16
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_16_opA.fifo),
        .read_port(rd_mul_18_16_opA.fifo)
        );        

        //line_buffer_0<->mul18_17
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_2_mul_18_17
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_17_opA.fifo),
        .read_port(rd_mul_18_17_opA.fifo)
        );

        //line_buffer_1<->mul18_18
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_2_mul_18_18
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_18_opA.fifo),
        .read_port(rd_mul_18_18_opA.fifo)
        );

        //line_buffer_2<->mul18_19
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_2_mul_18_19
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_19_opA.fifo),
        .read_port(rd_mul_18_19_opA.fifo)
        );

        //line_buffer_3<->mul18_20
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_2_mul_18_20
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_20_opA.fifo),
        .read_port(rd_mul_18_20_opA.fifo)
        );

        //line_buffer_4<->mul18_21
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_2_mul_18_21
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_21_opA.fifo),
        .read_port(rd_mul_18_21_opA.fifo)
        );

        //line_buffer_5<->mul18_22
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_2_mul_18_22
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_22_opA.fifo),
        .read_port(rd_mul_18_22_opA.fifo)
        );

        //line_buffer_6<->mul18_23
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_6_2_mul_18_23
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_line_buffer_6_2_out_pel.fifo),
        .read_port(rd_mul_18_23_opA.fifo)
        );

	//4� colonna
        
        //remove_h_3<->mul18_24
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_3_mul_18_24
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_24_opA.fifo),
        .read_port(rd_mul_18_24_opA.fifo)
        ); 

        //line_buffer_0<->mul18_25
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_3_mul_18_25
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_25_opA.fifo),
        .read_port(rd_mul_18_25_opA.fifo)
        );
        
        //line_buffer_1<->mul18_26
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_3_mul_18_26
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_26_opA.fifo),
        .read_port(rd_mul_18_26_opA.fifo)
        );

        //line_buffer_2<->mul18_27
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_3_mul_18_27
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_27_opA.fifo),
        .read_port(rd_mul_18_27_opA.fifo)
        );

        //line_buffer_3<->mul18_28
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_3_mul_18_28
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_28_opA.fifo),
        .read_port(rd_mul_18_28_opA.fifo)
        );

        
        //line_buffer_4<->mul18_29
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_3_mul_18_29
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_29_opA.fifo),
        .read_port(rd_mul_18_29_opA.fifo)
        );

        //line_buffer_5<->mul18_30
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_3_mul_18_30
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_30_opA.fifo),
        .read_port(rd_mul_18_30_opA.fifo)
        );

        //line_buffer_6<->mul18_31
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_6_3_mul_18_31
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_line_buffer_6_3_out_pel.fifo),
        .read_port(rd_mul_18_31_opA.fifo)
        );

    //5� colonna
    
        //remove_h4<->mul18_32
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_4_mul_18_32
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_32_opA.fifo),
        .read_port(rd_mul_18_32_opA.fifo)
        );

        //line_buffer_0<->mul18_33
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_4_mul_18_33
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_33_opA.fifo),
        .read_port(rd_mul_18_33_opA.fifo)
        );

        //line_buffer_1<->mul18_34
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_4_mul_18_34
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_34_opA.fifo),
        .read_port(rd_mul_18_34_opA.fifo)
        );

        //line_buffer_2<->mul18_35
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_4_mul_18_35
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_35_opA.fifo),
        .read_port(rd_mul_18_35_opA.fifo)
        );

        //line_buffer_3<->mul18_36
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_4_mul_18_36
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_36_opA.fifo),
        .read_port(rd_mul_18_36_opA.fifo)
        );

        //line_buffer_4<->mul18_37
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_4_mul_18_37
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_37_opA.fifo),
        .read_port(rd_mul_18_37_opA.fifo)
        );
		
        //line_buffer_5<->mul18_38
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_4_mul_18_38
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_38_opA.fifo),
        .read_port(rd_mul_18_38_opA.fifo)
        );		

        //line_buffer_6<->mul18_39
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_6_4_mul_18_39
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_line_buffer_6_4_out_pel.fifo),
        .read_port(rd_mul_18_39_opA.fifo)
        );

	//6� colonna

        //remove_h5<->mul18_40
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_5_mul_18_40
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_40_opA.fifo),
        .read_port(rd_mul_18_40_opA.fifo)
        );

        //line_buffer_0<->mul18_41
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_5_mul_18_41
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_41_opA.fifo),
        .read_port(rd_mul_18_41_opA.fifo)
        );

        //line_buffer_1<->mul18_42
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_5_mul_18_42
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_42_opA.fifo),
        .read_port(rd_mul_18_42_opA.fifo)
        );

        //line_buffer_2<->mul18_43
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_5_mul_18_43
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_43_opA.fifo),
        .read_port(rd_mul_18_43_opA.fifo)
        );

        //line_buffer_3<->mul18_44
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_5_mul_18_44
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_44_opA.fifo),
        .read_port(rd_mul_18_44_opA.fifo)
        );

        //line_buffer_4<->mul18_45
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_5_mul_18_45
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_45_opA.fifo),
        .read_port(rd_mul_18_45_opA.fifo)
        );
		
        //line_buffer_5<->mul18_46
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_5_mul_18_46
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_46_opA.fifo),
        .read_port(rd_mul_18_46_opA.fifo)
        );		

        //line_buffer_6<->mul18_47
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_6_5_mul_18_47
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_line_buffer_6_5_out_pel.fifo),
        .read_port(rd_mul_18_47_opA.fifo)
        );

	//7� colonna

        //remove6<->mul18_48
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_6_mul_18_48
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_48_opA.fifo),
        .read_port(rd_mul_18_48_opA.fifo)
        );
          
        //line_buffer_0<->mul18_49
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_6_mul_18_49
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_49_opA.fifo),
        .read_port(rd_mul_18_49_opA.fifo)
        );        

        //line_buffer_1<->mul18_50
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_6_mul_18_50
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_50_opA.fifo),
        .read_port(rd_mul_18_50_opA.fifo)
        );

        //line_buffer_2<->mul18_51
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_6_mul_18_51
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_51_opA.fifo),
        .read_port(rd_mul_18_51_opA.fifo)
        );
		
        //line_buffer_3<->mul18_52
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_6_mul_18_52
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_52_opA.fifo),
        .read_port(rd_mul_18_52_opA.fifo)
        );

        //line_buffer_4<->mul18_53
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_6_mul_18_53
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_53_opA.fifo),
        .read_port(rd_mul_18_53_opA.fifo)
        );		

        //line_buffer_5<->mul18_54
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_6_mul_18_54
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_54_opA.fifo),
        .read_port(rd_mul_18_54_opA.fifo)
        );

        //line_buffer_6<->mul18_55
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_6_6_mul_18_55
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_line_buffer_6_6_out_pel.fifo),
        .read_port(rd_mul_18_55_opA.fifo)
        );

    //8� colonna    
		
        //remove7<->mul18_56
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_7_mul_18_56
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_56_opA.fifo),
        .read_port(rd_mul_18_56_opA.fifo)
        );
            
         //line_buffer_0<->mul18_57
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_7_mul_18_57
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_57_opA.fifo),
        .read_port(rd_mul_18_57_opA.fifo)
        );          

       //line_buffer_1<->mul18_58
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_7_mul_18_58
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_58_opA.fifo),
        .read_port(rd_mul_18_58_opA.fifo)
        );   
                           
        //line_buffer_2<->mul18_59
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_7_mul_18_59
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_59_opA.fifo),
        .read_port(rd_mul_18_59_opA.fifo)
        );

        //line_buffer_3<->mul18_60
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_7_mul_18_60
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_60_opA.fifo),
        .read_port(rd_mul_18_60_opA.fifo)
        );

        //line_buffer_4<->mul18_61
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_7_mul_18_61
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_61_opA.fifo),
        .read_port(rd_mul_18_61_opA.fifo)
        );

        //line_buffer_5<->mul18_62
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_7_mul_18_62
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_62_opA.fifo),
        .read_port(rd_mul_18_62_opA.fifo)
        );

        //line_buffer_6<->mul18_63
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_6_7_mul_18_63
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_line_buffer_6_7_out_pel.fifo),
        .read_port(rd_mul_18_63_opA.fifo)
        );
        
   //coeff_v<->mul18 
    
    //1�riga 

        //coeff_luma_v<->mul_18_0
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_0_opB.fifo),
        .read_port(rd_mul_18_0_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_1
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_1_opB.fifo),
        .read_port(rd_mul_18_1_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_2
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_2_opB.fifo),
        .read_port(rd_mul_18_2_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_3
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_3_opB.fifo),
        .read_port(rd_mul_18_3_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_4
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_4_opB.fifo),
        .read_port(rd_mul_18_4_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_5
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_5_opB.fifo),
        .read_port(rd_mul_18_5_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_6
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_6_opB.fifo),
        .read_port(rd_mul_18_6_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_7
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_7_opB.fifo),
        .read_port(rd_mul_18_7_opB.fifo)
        );    
    
    //2� riga
    
        //coeff_luma_v<->mul_18_8
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_8
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_8_opB.fifo),
        .read_port(rd_mul_18_8_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_9
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_9
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_9_opB.fifo),
        .read_port(rd_mul_18_9_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_10
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_10
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_10_opB.fifo),
        .read_port(rd_mul_18_10_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_11
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_11
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_11_opB.fifo),
        .read_port(rd_mul_18_11_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_12
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_12
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_12_opB.fifo),
        .read_port(rd_mul_18_12_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_13
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_13
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_13_opB.fifo),
        .read_port(rd_mul_18_13_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_14
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_14
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_14_opB.fifo),
        .read_port(rd_mul_18_14_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_15
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_15
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_15_opB.fifo),
        .read_port(rd_mul_18_15_opB.fifo)
        );        
    
    //3� riga
    
        //coeff_luma_v<->mul_18_16
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_16
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_16_opB.fifo),
        .read_port(rd_mul_18_16_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_17
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_17
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_17_opB.fifo),
        .read_port(rd_mul_18_17_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_18
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_18
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_18_opB.fifo),
        .read_port(rd_mul_18_18_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_19
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_19
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_19_opB.fifo),
        .read_port(rd_mul_18_19_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_20
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_20
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_20_opB.fifo),
        .read_port(rd_mul_18_20_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_21
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_21
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_21_opB.fifo),
        .read_port(rd_mul_18_21_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_22
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_22
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_22_opB.fifo),
        .read_port(rd_mul_18_22_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_23
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_23
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_23_opB.fifo),
        .read_port(rd_mul_18_23_opB.fifo)
        );
            
    //4� riga
    
        //coeff_luma_v<->mul_18_24
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_24
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_24_opB.fifo),
        .read_port(rd_mul_18_24_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_25
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_25
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_25_opB.fifo),
        .read_port(rd_mul_18_25_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_26
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_26
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_26_opB.fifo),
        .read_port(rd_mul_18_26_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_27
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_27
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_27_opB.fifo),
        .read_port(rd_mul_18_27_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_28
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_28
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_28_opB.fifo),
        .read_port(rd_mul_18_28_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_29
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_29
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_29_opB.fifo),
        .read_port(rd_mul_18_29_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_30
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_30
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_30_opB.fifo),
        .read_port(rd_mul_18_30_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_31
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_31
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_31_opB.fifo),
        .read_port(rd_mul_18_31_opB.fifo)
        );
    
    //5� riga
    
        //coeff_luma_v<->mul_18_32
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_32
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_32_opB.fifo),
        .read_port(rd_mul_18_32_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_33
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_33
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_33_opB.fifo),
        .read_port(rd_mul_18_33_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_34
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_34
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_34_opB.fifo),
        .read_port(rd_mul_18_34_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_35
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_35
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_35_opB.fifo),
        .read_port(rd_mul_18_35_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_36
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_36
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_36_opB.fifo),
        .read_port(rd_mul_18_36_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_37
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_37
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_37_opB.fifo),
        .read_port(rd_mul_18_37_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_38
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_38
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_38_opB.fifo),
        .read_port(rd_mul_18_38_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_39
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_39
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_39_opB.fifo),
        .read_port(rd_mul_18_39_opB.fifo)
        );
    
    //6� riga
    
        //coeff_luma_v<->mul_18_40
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_40
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_40_opB.fifo),
        .read_port(rd_mul_18_40_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_41
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_41
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_41_opB.fifo),
        .read_port(rd_mul_18_41_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_42
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_42
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_42_opB.fifo),
        .read_port(rd_mul_18_42_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_43
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_43
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_43_opB.fifo),
        .read_port(rd_mul_18_43_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_44
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_44
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_44_opB.fifo),
        .read_port(rd_mul_18_44_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_45
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_45
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_45_opB.fifo),
        .read_port(rd_mul_18_45_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_46
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_46
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_46_opB.fifo),
        .read_port(rd_mul_18_46_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_47
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_47
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_47_opB.fifo),
        .read_port(rd_mul_18_47_opB.fifo)
        );
        
    //7� riga
    
        //coeff_luma_v<->mul_18_48
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_48
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_48_opB.fifo),
        .read_port(rd_mul_18_48_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_49
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_49
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_49_opB.fifo),
        .read_port(rd_mul_18_49_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_50
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_50
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_50_opB.fifo),
        .read_port(rd_mul_18_50_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_51
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_51
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_51_opB.fifo),
        .read_port(rd_mul_18_51_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_52
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_52
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_52_opB.fifo),
        .read_port(rd_mul_18_52_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_53
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_53
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_53_opB.fifo),
        .read_port(rd_mul_18_53_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_54
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_54
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_54_opB.fifo),
        .read_port(rd_mul_18_54_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_55
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_55
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_55_opB.fifo),
        .read_port(rd_mul_18_55_opB.fifo)
        );
            
    //8�riga
        
        //coeff_luma_v<->mul_18_56
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_56
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_56_opB.fifo),
        .read_port(rd_mul_18_56_opB.fifo)
        );        
        
        //coeff_luma_v<->mul_18_57
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_57
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_57_opB.fifo),
        .read_port(rd_mul_18_57_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_58
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_58
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_58_opB.fifo),
        .read_port(rd_mul_18_58_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_59
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_59
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_59_opB.fifo),
        .read_port(rd_mul_18_59_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_60
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_60
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_60_opB.fifo),
        .read_port(rd_mul_18_60_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_61
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_61
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_61_opB.fifo),
        .read_port(rd_mul_18_61_opB.fifo)
        );
        
        //coeff_luma_v<->mul_18_62
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_62
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_62_opB.fifo),
        .read_port(rd_mul_18_62_opB.fifo)
        );        

        //coeff_luma_v<->mul_18_63
        fifo_ms #(9,DEPTH,FLUX) fifo_coeff_luma_v_mul_18_63
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_mul_18_63_opB.fifo),
        .read_port(rd_mul_18_63_opB.fifo)
        );        

    //LIME: INPUT REALSIZE LINE BUFFER (x7)
        
        //derive_real_size<->line_buffer_0
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_line_buffer_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_0_real_size.fifo),
        .read_port(rd_line_buffer_0_real_size.fifo)
        );

        //derive_real_size<->line_buffer_1
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_line_buffer_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_1_real_size.fifo),
        .read_port(rd_line_buffer_1_real_size.fifo)
        );
        
        //derive_real_size<->line_buffer_2
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_line_buffer_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_2_real_size.fifo),
        .read_port(rd_line_buffer_2_real_size.fifo)
        );

        //derive_real_size<->line_buffer_3
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_line_buffer_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_3_real_size.fifo),
        .read_port(rd_line_buffer_3_real_size.fifo)
        );  
        //derive_real_size<->line_buffer_4
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_line_buffer_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_4_real_size.fifo),
        .read_port(rd_line_buffer_4_real_size.fifo)
        );

        //derive_real_size<->line_buffer_5
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_line_buffer_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_5_real_size.fifo),
        .read_port(rd_line_buffer_5_real_size.fifo)
        );
        
        //derive_real_size<->line_buffer_6
        fifo_ms #(7,DEPTH,FLUX) fifo_derive_real_size_line_buffer_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_6_real_size.fifo),
        .read_port(rd_line_buffer_6_real_size.fifo)
        );        
                
    //LIGHT BLUE: INPUT EXTSIZE LINE BUFFER (x7)
        
        //extsize<->line_buffer_0
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_linebuffer0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_0_ext_size.fifo),
        .read_port(rd_line_buffer_0_ext_size.fifo)
        );    

        //extsize<->line_buffer_1
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_linebuffer1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_1_ext_size.fifo),
        .read_port(rd_line_buffer_1_ext_size.fifo)
        );

        //extsize<->line_buffer_2
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_linebuffer2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_2_ext_size.fifo),
        .read_port(rd_line_buffer_2_ext_size.fifo)
        );

        //extsize<->line_buffer_3
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_linebuffer3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_3_ext_size.fifo),
        .read_port(rd_line_buffer_3_ext_size.fifo)
        );

        //extsize<->line_buffer_4
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_linebuffer4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_4_ext_size.fifo),
        .read_port(rd_line_buffer_4_ext_size.fifo)
        );

        //extsize<->line_buffer_5
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_linebuffer5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_5_ext_size.fifo),
        .read_port(rd_line_buffer_5_ext_size.fifo)
        );

        //extsize<->line_buffer_6
        fifo_ms #(7,DEPTH,FLUX) fifo_extsize_linebuffer6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_6_ext_size.fifo),
        .read_port(rd_line_buffer_6_ext_size.fifo)
        );
		
	//remove_h<->line_buffer_0
		
       //remove_h_0<->line_buffer_0_0
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_0_line_buffer_0_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_0_0_in_pel.fifo),
        .read_port(rd_line_buffer_0_0_in_pel.fifo)
        );    

       //remove_h_1<->line_buffer_0_1
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_1_line_buffer_0_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_0_1_in_pel.fifo),
        .read_port(rd_line_buffer_0_1_in_pel.fifo)
        );    

       //remove_h_2<->line_buffer_0_2
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_2_line_buffer_0_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_0_2_in_pel.fifo),
        .read_port(rd_line_buffer_0_2_in_pel.fifo)
        );    

       //remove_h_3<->line_buffer_0_3
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_3_line_buffer_0_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_0_3_in_pel.fifo),
        .read_port(rd_line_buffer_0_3_in_pel.fifo)
        );    

       //remove_h_4<->line_buffer_0_4
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_4_line_buffer_0_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_0_4_in_pel.fifo),
        .read_port(rd_line_buffer_0_4_in_pel.fifo)
        );    
		
       //remove_h_5<->line_buffer_0_5
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_5_line_buffer_0_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_0_5_in_pel.fifo),
        .read_port(rd_line_buffer_0_5_in_pel.fifo)
        );    

       //remove_h_6<->line_buffer_0_6
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_6_line_buffer_0_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_0_6_in_pel.fifo),
        .read_port(rd_line_buffer_0_6_in_pel.fifo)
        );    		

       //remove_h_7<->line_buffer_0_7
        fifo_ms #(18,DEPTH,FLUX) fifo_remove_h_7_line_buffer_0_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_0_7_in_pel.fifo),
        .read_port(rd_line_buffer_0_7_in_pel.fifo)
        );    


	//line_buffer_0<->line_buffer_1
		
       //line_buffer_0_0<->line_buffer_1_0
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_0_line_buffer_1_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_1_0_in_pel.fifo),
        .read_port(rd_line_buffer_1_0_in_pel.fifo)
        );    

       //line_buffer_0_1<->line_buffer_1_1
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_1_line_buffer_1_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_1_1_in_pel.fifo),
        .read_port(rd_line_buffer_1_1_in_pel.fifo)
        );    

       //line_buffer_0_2<->line_buffer_1_2
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_2_line_buffer_1_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_1_2_in_pel.fifo),
        .read_port(rd_line_buffer_1_2_in_pel.fifo)
        );    

       //line_buffer_0_3<->line_buffer_1_3
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_3_line_buffer_1_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_1_3_in_pel.fifo),
        .read_port(rd_line_buffer_1_3_in_pel.fifo)
        );    

       //line_buffer_0_4<->line_buffer_1_4
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_4_line_buffer_1_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_1_4_in_pel.fifo),
        .read_port(rd_line_buffer_1_4_in_pel.fifo)
        );    
		
       //line_buffer_0_5<->line_buffer_1_5
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_5_line_buffer_1_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_1_5_in_pel.fifo),
        .read_port(rd_line_buffer_1_5_in_pel.fifo)
        );    

       //line_buffer_0_6<->line_buffer_1_6
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_6_line_buffer_1_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_1_6_in_pel.fifo),
        .read_port(rd_line_buffer_1_6_in_pel.fifo)
        );    		

       //line_buffer_0_7<->line_buffer_1_7
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_0_7_line_buffer_1_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_1_7_in_pel.fifo),
        .read_port(rd_line_buffer_1_7_in_pel.fifo)
        );    


	//line_buffer_1<->line_buffer_2
		
       //line_buffer_1_0<->line_buffer_2_0
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_0_line_buffer_2_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_2_0_in_pel.fifo),
        .read_port(rd_line_buffer_2_0_in_pel.fifo)
        );    

       //line_buffer_1_1<->line_buffer_2_1
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_1_line_buffer_2_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_2_1_in_pel.fifo),
        .read_port(rd_line_buffer_2_1_in_pel.fifo)
        );    

       //line_buffer_1_2<->line_buffer_2_2
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_2_line_buffer_2_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_2_2_in_pel.fifo),
        .read_port(rd_line_buffer_2_2_in_pel.fifo)
        );    

       //line_buffer_1_3<->line_buffer_2_3
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_3_line_buffer_2_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_2_3_in_pel.fifo),
        .read_port(rd_line_buffer_2_3_in_pel.fifo)
        );    

       //line_buffer_1_4<->line_buffer_2_4
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_4_line_buffer_2_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_2_4_in_pel.fifo),
        .read_port(rd_line_buffer_2_4_in_pel.fifo)
        );    
		
       //line_buffer_1_5<->line_buffer_2_5
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_5_line_buffer_2_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_2_5_in_pel.fifo),
        .read_port(rd_line_buffer_2_5_in_pel.fifo)
        );    

       //line_buffer_1_6<->line_buffer_2_6
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_6_line_buffer_2_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_2_6_in_pel.fifo),
        .read_port(rd_line_buffer_2_6_in_pel.fifo)
        );    		

       //line_buffer_1_7<->line_buffer_2_7
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_1_7_line_buffer_2_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_2_7_in_pel.fifo),
        .read_port(rd_line_buffer_2_7_in_pel.fifo)
        );



	//line_buffer_2<->line_buffer_3
		
       //line_buffer_2_0<->line_buffer_3_0
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_0_line_buffer_3_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_3_0_in_pel.fifo),
        .read_port(rd_line_buffer_3_0_in_pel.fifo)
        );    

       //line_buffer_2_1<->line_buffer_3_1
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_1_line_buffer_3_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_3_1_in_pel.fifo),
        .read_port(rd_line_buffer_3_1_in_pel.fifo)
        );    

       //line_buffer_2_2<->line_buffer_3_2
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_2_line_buffer_3_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_3_2_in_pel.fifo),
        .read_port(rd_line_buffer_3_2_in_pel.fifo)
        );    

       //line_buffer_2_3<->line_buffer_3_3
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_3_line_buffer_3_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_3_3_in_pel.fifo),
        .read_port(rd_line_buffer_3_3_in_pel.fifo)
        );    

       //line_buffer_2_4<->line_buffer_3_4
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_4_line_buffer_3_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_3_4_in_pel.fifo),
        .read_port(rd_line_buffer_3_4_in_pel.fifo)
        );    
		
       //line_buffer_2_5<->line_buffer_3_5
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_5_line_buffer_3_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_3_5_in_pel.fifo),
        .read_port(rd_line_buffer_3_5_in_pel.fifo)
        );    

       //line_buffer_2_6<->line_buffer_3_6
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_6_line_buffer_3_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_3_6_in_pel.fifo),
        .read_port(rd_line_buffer_3_6_in_pel.fifo)
        );    		

       //line_buffer_2_7<->line_buffer_3_7
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_2_7_line_buffer_3_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_3_7_in_pel.fifo),
        .read_port(rd_line_buffer_3_7_in_pel.fifo)
        );



	//line_buffer_3<->line_buffer_4
		
       //line_buffer_3_0<->line_buffer_4_0
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_0_line_buffer_4_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_4_0_in_pel.fifo),
        .read_port(rd_line_buffer_4_0_in_pel.fifo)
        );    

       //line_buffer_3_1<->line_buffer_4_1
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_1_line_buffer_4_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_4_1_in_pel.fifo),
        .read_port(rd_line_buffer_4_1_in_pel.fifo)
        );    

       //line_buffer_3_2<->line_buffer_4_2
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_2_line_buffer_4_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_4_2_in_pel.fifo),
        .read_port(rd_line_buffer_4_2_in_pel.fifo)
        );    

       //line_buffer_3_3<->line_buffer_4_3
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_3_line_buffer_4_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_4_3_in_pel.fifo),
        .read_port(rd_line_buffer_4_3_in_pel.fifo)
        );    

       //line_buffer_3_4<->line_buffer_4_4
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_4_line_buffer_4_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_4_4_in_pel.fifo),
        .read_port(rd_line_buffer_4_4_in_pel.fifo)
        );    
		
       //line_buffer_3_5<->line_buffer_4_5
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_5_line_buffer_4_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_4_5_in_pel.fifo),
        .read_port(rd_line_buffer_4_5_in_pel.fifo)
        );    

       //line_buffer_3_6<->line_buffer_4_6
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_6_line_buffer_4_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_4_6_in_pel.fifo),
        .read_port(rd_line_buffer_4_6_in_pel.fifo)
        );    		

       //line_buffer_3_7<->line_buffer_4_7
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_3_7_line_buffer_4_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_4_7_in_pel.fifo),
        .read_port(rd_line_buffer_4_7_in_pel.fifo)
        );
		
		

	//line_buffer_4<->line_buffer_5
		
       //line_buffer_4_0<->line_buffer_5_0
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_0_line_buffer_5_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_5_0_in_pel.fifo),
        .read_port(rd_line_buffer_5_0_in_pel.fifo)
        );    

       //line_buffer_4_1<->line_buffer_5_1
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_1_line_buffer_5_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_5_1_in_pel.fifo),
        .read_port(rd_line_buffer_5_1_in_pel.fifo)
        );    

       //line_buffer_4_2<->line_buffer_5_2
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_2_line_buffer_5_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_5_2_in_pel.fifo),
        .read_port(rd_line_buffer_5_2_in_pel.fifo)
        );    

       //line_buffer_4_3<->line_buffer_5_3
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_3_line_buffer_5_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_5_3_in_pel.fifo),
        .read_port(rd_line_buffer_5_3_in_pel.fifo)
        );    

       //line_buffer_4_4<->line_buffer_5_4
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_4_line_buffer_5_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_5_4_in_pel.fifo),
        .read_port(rd_line_buffer_5_4_in_pel.fifo)
        );    
		
       //line_buffer_4_5<->line_buffer_5_5
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_5_line_buffer_5_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_5_5_in_pel.fifo),
        .read_port(rd_line_buffer_5_5_in_pel.fifo)
        );    

       //line_buffer_4_6<->line_buffer_5_6
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_6_line_buffer_5_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_5_6_in_pel.fifo),
        .read_port(rd_line_buffer_5_6_in_pel.fifo)
        );    		

       //line_buffer_4_7<->line_buffer_5_7
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_4_7_line_buffer_5_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_5_7_in_pel.fifo),
        .read_port(rd_line_buffer_5_7_in_pel.fifo)
        );		
		
		

	//line_buffer_5<->line_buffer_6
		
       //line_buffer_5_0<->line_buffer_6_0
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_0_line_buffer_6_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_6_0_in_pel.fifo),
        .read_port(rd_line_buffer_6_0_in_pel.fifo)
        );    

       //line_buffer_5_1<->line_buffer_6_1
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_1_line_buffer_6_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_6_1_in_pel.fifo),
        .read_port(rd_line_buffer_6_1_in_pel.fifo)
        );    

       //line_buffer_5_2<->line_buffer_6_2
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_2_line_buffer_6_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_6_2_in_pel.fifo),
        .read_port(rd_line_buffer_6_2_in_pel.fifo)
        );    

       //line_buffer_5_3<->line_buffer_6_3
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_3_line_buffer_6_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_6_3_in_pel.fifo),
        .read_port(rd_line_buffer_6_3_in_pel.fifo)
        );    

       //line_buffer_5_4<->line_buffer_6_4
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_4_line_buffer_6_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_6_4_in_pel.fifo),
        .read_port(rd_line_buffer_6_4_in_pel.fifo)
        );    
		
       //line_buffer_5_5<->line_buffer_6_5
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_5_line_buffer_6_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_6_5_in_pel.fifo),
        .read_port(rd_line_buffer_6_5_in_pel.fifo)
        );    

       //line_buffer_5_6<->line_buffer_6_6
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_6_line_buffer_6_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_6_6_in_pel.fifo),
        .read_port(rd_line_buffer_6_6_in_pel.fifo)
        );    		

       //line_buffer_5_7<->line_buffer_6_7
        fifo_ms #(18,DEPTH,FLUX) fifo_line_buffer_5_7_line_buffer_6_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_fifo_line_buffer_6_7_in_pel.fifo),
        .read_port(rd_line_buffer_6_7_in_pel.fifo)
        );

        
    //1� adder tree
        //mul_18_0<->adder_27_0
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_0_add_27_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_0_prod.fifo),
        .read_port(rd_add_27_0_opA.fifo)
        );

        //mul_18_1<->adder_27_0
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_1_add_27_0
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_1_prod.fifo),
        .read_port(rd_add_27_0_opB.fifo)
        );
        
        //mul_18_2<->adder_27_1
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_2_add_27_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_2_prod.fifo),
        .read_port(rd_add_27_1_opA.fifo)
        );  

        //mul_18_3<->adder_27_1
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_3_add_27_1
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_3_prod.fifo),
        .read_port(rd_add_27_1_opB.fifo)
        );

        //mul_18_4<->adder_27_2
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_4_add_27_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_4_prod.fifo),
        .read_port(rd_add_27_2_opA.fifo)
        );
        
        //mul_18_5<->adder_27_2
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_5_add_27_2
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_5_prod.fifo),
        .read_port(rd_add_27_2_opB.fifo)
        );

        //mul_18_6<->adder_27_3
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_6_add_27_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_6_prod.fifo),
        .read_port(rd_add_27_3_opA.fifo)
        );
        
        //mul_18_7<->adder_27_3
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_7_add_27_3
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_7_prod.fifo),
        .read_port(rd_add_27_3_opB.fifo)
        );

        //adder_27_0<->adder_27_4
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_0_add_27_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_0_sum.fifo),
        .read_port(rd_add_27_4_opA.fifo)
        );  

        //adder_27_1<->adder_27_4
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_1_add_27_4
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_1_sum.fifo),
        .read_port(rd_add_27_4_opB.fifo)
        );

        //adder_27_2<->adder_27_5
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_2_add_27_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_2_sum.fifo),
        .read_port(rd_add_27_5_opA.fifo)
        );
        
        //adder_27_3<->adder_27_5
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_3_add_27_5
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_3_sum.fifo),
        .read_port(rd_add_27_5_opB.fifo)
        );

        //adder_27_4<->adder_27_6
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_4_add_27_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_4_sum.fifo),
        .read_port(rd_add_27_6_opA.fifo)
        );
        
        //adder_27_5<->adder_27_6
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_5_add_27_6
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_5_sum.fifo),
        .read_port(rd_add_27_6_opB.fifo)
        );

    
    //2� adder tree

        //mul_18_8<->adder_27_7
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_8_add_27_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_8_prod.fifo),
        .read_port(rd_add_27_7_opA.fifo)
        );

        //mul_18_9<->adder_27_7
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_9_add_27_7
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_9_prod.fifo),
        .read_port(rd_add_27_7_opB.fifo)
        );
        
        //mul_18_10<->adder_27_8
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_10_9_add_27_8
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_10_prod.fifo),
        .read_port(rd_add_27_8_opA.fifo)
        );  

        //mul_18_11<->adder_27_8
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_11_add_27_8
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_11_prod.fifo),
        .read_port(rd_add_27_8_opB.fifo)
        );

        //mul_18_12<->adder_27_9
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_12_add_27_9
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_12_prod.fifo),
        .read_port(rd_add_27_9_opA.fifo)
        );
        
        //mul_18_13<->adder_27_9
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_13_add_27_9
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_13_prod.fifo),
        .read_port(rd_add_27_9_opB.fifo)
        );

        //mul_18_14<->adder_27_10
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_14_add_27_10
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_14_prod.fifo),
        .read_port(rd_add_27_10_opA.fifo)
        );
        
        //mul_18_15<->adder_27_10
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_15_add_27_10
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_15_prod.fifo),
        .read_port(rd_add_27_10_opB.fifo)
        );

        //adder_27_7<->adder_27_11
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_7_add_27_11
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_7_sum.fifo),
        .read_port(rd_add_27_11_opA.fifo)
        );  

        //adder_27_8<->adder_27_11
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_8_add_27_11
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_8_sum.fifo),
        .read_port(rd_add_27_11_opB.fifo)
        );

        //adder_27_9<->adder_27_12
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_9_add_27_12
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_9_sum.fifo),
        .read_port(rd_add_27_12_opA.fifo)
        );
        
        //adder_27_10<->adder_27_12
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_10_add_27_12
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_10_sum.fifo),
        .read_port(rd_add_27_12_opB.fifo)
        );

        //adder_27_11<->adder_27_13
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_11_add_27_13
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_11_sum.fifo),
        .read_port(rd_add_27_13_opA.fifo)
        );
        
        //adder_27_12<->adder_27_13
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_12_add_27_13
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_12_sum.fifo),
        .read_port(rd_add_27_13_opB.fifo)
        );
    
    //3� adder tree

        //mul_18_16<->adder_27_14
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_16_add_27_14
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_16_prod.fifo),
        .read_port(rd_add_27_14_opA.fifo)
        );

        //mul_18_17<->adder_27_14
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_17_add_27_14
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_17_prod.fifo),
        .read_port(rd_add_27_14_opB.fifo)
        );
        
        //mul_18_18<->adder_27_15
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_18_add_27_15
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_18_prod.fifo),
        .read_port(rd_add_27_15_opA.fifo)
        );  

        //mul_18_19<->adder_27_15
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_19_add_27_15
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_19_prod.fifo),
        .read_port(rd_add_27_15_opB.fifo)
        );

        //mul_18_20<->adder_27_16
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_20_add_27_16
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_20_prod.fifo),
        .read_port(rd_add_27_16_opA.fifo)
        );
        
        //mul_18_21<->adder_27_16
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_21_add_27_16
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_21_prod.fifo),
        .read_port(rd_add_27_16_opB.fifo)
        );

        //mul_18_22<->adder_27_17
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_22_add_27_17
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_22_prod.fifo),
        .read_port(rd_add_27_17_opA.fifo)
        );
        
        //mul_18_23<->adder_27_17
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_23_add_27_17
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_23_prod.fifo),
        .read_port(rd_add_27_17_opB.fifo)
        );

        //adder_27_14<->adder_27_18
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_14_add_27_18
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_14_sum.fifo),
        .read_port(rd_add_27_18_opA.fifo)
        );  

        //adder_27_15<->adder_27_18
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_15_add_27_18
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_15_sum.fifo),
        .read_port(rd_add_27_18_opB.fifo)
        );

        //adder_27_16<->adder_27_19
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_16_add_27_19
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_16_sum.fifo),
        .read_port(rd_add_27_19_opA.fifo)
        );
        
        //adder_27_17<->adder_27_19
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_17_add_27_19
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_17_sum.fifo),
        .read_port(rd_add_27_19_opB.fifo)
        );

        //adder_27_18<->adder_27_20
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_18_add_27_20
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_18_sum.fifo),
        .read_port(rd_add_27_20_opA.fifo)
        );
        
        //adder_27_19<->adder_27_20
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_19_add_27_20
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_19_sum.fifo),
        .read_port(rd_add_27_20_opB.fifo)
        );

    
    //4� adder tree

        //mul_18_24<->adder_27_21
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_24_add_27_21
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_24_prod.fifo),
        .read_port(rd_add_27_21_opA.fifo)
        );

        //mul_18_25<->adder_27_21
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_25_add_27_21
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_25_prod.fifo),
        .read_port(rd_add_27_21_opB.fifo)
        );
        
        //mul_18_26<->adder_27_22
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_26_add_27_22
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_26_prod.fifo),
        .read_port(rd_add_27_22_opA.fifo)
        );  

        //mul_18_27<->adder_27_22
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_27_add_27_22
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_27_prod.fifo),
        .read_port(rd_add_27_22_opB.fifo)
        );

        //mul_18_28<->adder_27_23
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_28_add_27_23
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_28_prod.fifo),
        .read_port(rd_add_27_23_opA.fifo)
        );
        
        //mul_18_29<->adder_27_23
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_29_add_27_23
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_29_prod.fifo),
        .read_port(rd_add_27_23_opB.fifo)
        );

        //mul_18_30<->adder_27_24
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_30_add_27_24
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_30_prod.fifo),
        .read_port(rd_add_27_24_opA.fifo)
        );
        
        //mul_18_31<->adder_27_24
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_31_add_27_24
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_31_prod.fifo),
        .read_port(rd_add_27_24_opB.fifo)
        );

        //adder_27_21<->adder_27_25
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_21_add_27_25
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_21_sum.fifo),
        .read_port(rd_add_27_25_opA.fifo)
        );  

        //adder_27_22<->adder_27_25
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_22_add_27_25
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_22_sum.fifo),
        .read_port(rd_add_27_25_opB.fifo)
        );

        //adder_27_23<->adder_27_26
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_23_add_27_26
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_23_sum.fifo),
        .read_port(rd_add_27_26_opA.fifo)
        );
        
        //adder_27_24<->adder_27_26
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_24_add_27_26
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_24_sum.fifo),
        .read_port(rd_add_27_26_opB.fifo)
        );

        //adder_27_25<->adder_27_27
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_25_add_27_27
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_25_sum.fifo),
        .read_port(rd_add_27_27_opA.fifo)
        );
        
        //adder_27_26<->adder_27_27
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_26_add_27_27
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_26_sum.fifo),
        .read_port(rd_add_27_27_opB.fifo)
        );
    
    //5� adder tree

        //mul_18_32<->adder_27_28
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_32_add_27_28
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_32_prod.fifo),
        .read_port(rd_add_27_28_opA.fifo)
        );

        //mul_18_33<->adder_27_28
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_33_add_27_28
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_33_prod.fifo),
        .read_port(rd_add_27_28_opB.fifo)
        );
        
        //mul_18_34<->adder_27_29
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_34_add_27_29
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_34_prod.fifo),
        .read_port(rd_add_27_29_opA.fifo)
        );  

        //mul_18_35<->adder_27_29
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_35_add_27_29
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_35_prod.fifo),
        .read_port(rd_add_27_29_opB.fifo)
        );

        //mul_18_36<->adder_27_30
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_36_add_27_30
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_36_prod.fifo),
        .read_port(rd_add_27_30_opA.fifo)
        );
        
        //mul_18_37<->adder_27_30
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_37_add_27_30
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_37_prod.fifo),
        .read_port(rd_add_27_30_opB.fifo)
        );

        //mul_18_38<->adder_27_31
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_38_add_27_31
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_38_prod.fifo),
        .read_port(rd_add_27_31_opA.fifo)
        );
        
        //mul_18_39<->adder_27_31
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_39_add_27_31
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_39_prod.fifo),
        .read_port(rd_add_27_31_opB.fifo)
        );

        //adder_27_28<->adder_27_32
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_28_add_27_32
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_28_sum.fifo),
        .read_port(rd_add_27_32_opA.fifo)
        );  

        //adder_27_29<->adder_27_32
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_29_add_27_32
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_29_sum.fifo),
        .read_port(rd_add_27_32_opB.fifo)
        );

        //adder_27_30<->adder_27_33
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_30_add_27_33
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_30_sum.fifo),
        .read_port(rd_add_27_33_opA.fifo)
        );
        
        //adder_27_31<->adder_27_33
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_31_add_27_33
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_31_sum.fifo),
        .read_port(rd_add_27_33_opB.fifo)
        );

        //adder_27_32<->adder_27_34
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_32_add_27_34
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_32_sum.fifo),
        .read_port(rd_add_27_34_opA.fifo)
        );
        
        //adder_27_33<->adder_27_34
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_33_add_27_34
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_33_sum.fifo),
        .read_port(rd_add_27_34_opB.fifo)
        );
    
    //6� adder tree

        //mul_18_40<->adder_27_35
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_40_add_27_35
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_40_prod.fifo),
        .read_port(rd_add_27_35_opA.fifo)
        );

        //mul_18_41<->adder_27_35
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_41_add_27_35
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_41_prod.fifo),
        .read_port(rd_add_27_35_opB.fifo)
        );
        
        //mul_18_42<->adder_27_36
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_42_add_27_36
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_42_prod.fifo),
        .read_port(rd_add_27_36_opA.fifo)
        );  

        //mul_18_43<->adder_27_36
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_43_add_27_36
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_43_prod.fifo),
        .read_port(rd_add_27_36_opB.fifo)
        );

        //mul_18_44<->adder_27_37
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_44_add_27_37
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_44_prod.fifo),
        .read_port(rd_add_27_37_opA.fifo)
        );
        
        //mul_18_45<->adder_27_37
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_45_add_27_37
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_45_prod.fifo),
        .read_port(rd_add_27_37_opB.fifo)
        );

        //mul_18_46<->adder_27_38
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_46_add_27_38
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_46_prod.fifo),
        .read_port(rd_add_27_38_opA.fifo)
        );
        
        //mul_18_47<->adder_27_38
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_47_add_27_38
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_47_prod.fifo),
        .read_port(rd_add_27_38_opB.fifo)
        );

        //adder_27_35<->adder_27_39
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_35_add_27_39
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_35_sum.fifo),
        .read_port(rd_add_27_39_opA.fifo)
        );  

        //adder_27_36<->adder_27_39
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_36_add_27_39
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_36_sum.fifo),
        .read_port(rd_add_27_39_opB.fifo)
        );

        //adder_27_37<->adder_27_40
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_37_add_27_40
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_37_sum.fifo),
        .read_port(rd_add_27_40_opA.fifo)
        );
        
        //adder_27_38<->adder_27_40
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_38_add_27_40
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_38_sum.fifo),
        .read_port(rd_add_27_40_opB.fifo)
        );

        //adder_27_39<->adder_27_41
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_39_add_27_41
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_39_sum.fifo),
        .read_port(rd_add_27_41_opA.fifo)
        );
        
        //adder_27_40<->adder_27_41
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_40_add_27_41
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_40_sum.fifo),
        .read_port(rd_add_27_41_opB.fifo)
        );
    
    //7� adder tree

        //mul_18_48<->adder_27_42
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_48_add_27_42
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_48_prod.fifo),
        .read_port(rd_add_27_42_opA.fifo)
        );

        //mul_18_49<->adder_27_42
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_49_add_27_42
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_49_prod.fifo),
        .read_port(rd_add_27_42_opB.fifo)
        );
        
        //mul_18_50<->adder_27_43
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_50_add_27_43
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_50_prod.fifo),
        .read_port(rd_add_27_43_opA.fifo)
        );  

        //mul_18_51<->adder_27_43
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_51_add_27_43
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_51_prod.fifo),
        .read_port(rd_add_27_43_opB.fifo)
        );

        //mul_18_52<->adder_27_44
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_52_add_27_44
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_52_prod.fifo),
        .read_port(rd_add_27_44_opA.fifo)
        );
        
        //mul_18_53<->adder_27_44
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_53_add_27_44
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_53_prod.fifo),
        .read_port(rd_add_27_44_opB.fifo)
        );

        //mul_18_54<->adder_27_45
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_54_add_27_45
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_54_prod.fifo),
        .read_port(rd_add_27_45_opA.fifo)
        );
        
        //mul_18_55<->adder_27_45
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_55_add_27_45
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_55_prod.fifo),
        .read_port(rd_add_27_45_opB.fifo)
        );

        //adder_27_42<->adder_27_46
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_42_add_27_46
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_42_sum.fifo),
        .read_port(rd_add_27_46_opA.fifo)
        );  

        //adder_27_43<->adder_27_46
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_43_add_27_46
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_43_sum.fifo),
        .read_port(rd_add_27_46_opB.fifo)
        );

        //adder_27_44<->adder_27_47
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_44_add_27_47
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_44_sum.fifo),
        .read_port(rd_add_27_47_opA.fifo)
        );
        
        //adder_27_45<->adder_27_47
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_45_add_27_47
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_45_sum.fifo),
        .read_port(rd_add_27_47_opB.fifo)
        );

        //adder_27_46<->adder_27_48
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_46_add_27_48
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_46_sum.fifo),
        .read_port(rd_add_27_48_opA.fifo)
        );
        
        //adder_27_47<->adder_27_48
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_47_add_27_48
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_47_sum.fifo),
        .read_port(rd_add_27_48_opB.fifo)
        );
    
    //8� adder tree       

        //mul_18_56<->adder_27_49
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_56_add_27_49
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_56_prod.fifo),
        .read_port(rd_add_27_49_opA.fifo)
        );

        //mul_18_57<->adder_27_49
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_57_add_27_49
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_57_prod.fifo),
        .read_port(rd_add_27_49_opB.fifo)
        );
        
        //mul_18_58<->adder_27_50
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_58_add_27_50
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_58_prod.fifo),
        .read_port(rd_add_27_50_opA.fifo)
        );  

        //mul_18_59<->adder_27_50
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_59_add_27_50
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_59_prod.fifo),
        .read_port(rd_add_27_50_opB.fifo)
        );

        //mul_18_60<->adder_27_51
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_60_add_27_51
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_60_prod.fifo),
        .read_port(rd_add_27_51_opA.fifo)
        );
        
        //mul_18_61<->adder_27_51
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_61_add_27_51
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_61_prod.fifo),
        .read_port(rd_add_27_51_opB.fifo)
        );

        //mul_18_62<->adder_27_52
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_62_add_27_52
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_62_prod.fifo),
        .read_port(rd_add_27_52_opA.fifo)
        );
        
        //mul_18_63<->adder_27_52
        fifo_ms #(27,DEPTH,FLUX) fifo_mul_18_63_add_27_52
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_mul_18_63_prod.fifo),
        .read_port(rd_add_27_52_opB.fifo)
        );

        //adder_27_49<->adder_27_53
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_49_add_27_53
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_49_sum.fifo),
        .read_port(rd_add_27_53_opA.fifo)
        );  

        //adder_27_50<->adder_27_53
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_50_add_27_53
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_50_sum.fifo),
        .read_port(rd_add_27_53_opB.fifo)
        );

        //adder_27_51<->adder_27_54
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_51_add_27_54
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_51_sum.fifo),
        .read_port(rd_add_27_54_opA.fifo)
        );
        
        //adder_27_52<->adder_27_54
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_52_add_27_54
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_52_sum.fifo),
        .read_port(rd_add_27_54_opB.fifo)
        );

        //adder_27_53<->adder_27_55
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_53_add_27_55
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_53_sum.fifo),
        .read_port(rd_add_27_55_opA.fifo)
        );
        
        //adder_27_54<->adder_27_55
        fifo_ms #(27,DEPTH,FLUX) fifo_add_27_54_add_27_55
        (
        .clk(clk),
        .rst(rst),
        .write_port(wr_add_27_54_sum.fifo),
        .read_port(rd_add_27_55_opB.fifo)
        );



//FINE FIFO SECONDA PARTE




//MODULI SECONDA PARTE



       //LINE BUFFER (x7); I: LIME (1�HALF) / LIGHT BLUE (1�HALF) / RED (1�-2�HALF) - O: DARK GREY / RED

        //line_buffer_0
        line_buffer_8p#(FLUX) line_buffer0
        (
        .clk(clk),
        .rst(rst),        
        .read_port_real_size(rd_line_buffer_0_real_size.actor),
        .read_port_ext_size(rd_line_buffer_0_ext_size.actor),
        .read_port_in_pel_0(rd_line_buffer_0_0_in_pel.actor),            
		.read_port_in_pel_1(rd_line_buffer_0_1_in_pel.actor),            
		.read_port_in_pel_2(rd_line_buffer_0_2_in_pel.actor),            
		.read_port_in_pel_3(rd_line_buffer_0_3_in_pel.actor),            
		.read_port_in_pel_4(rd_line_buffer_0_4_in_pel.actor),            
		.read_port_in_pel_5(rd_line_buffer_0_5_in_pel.actor),            
		.read_port_in_pel_6(rd_line_buffer_0_6_in_pel.actor),            
		.read_port_in_pel_7(rd_line_buffer_0_7_in_pel.actor),
		.write_port_out_pel_0(wr_line_buffer_0_0_out_pel.actor),        		
        .write_port_out_pel_1(wr_line_buffer_0_1_out_pel.actor),        
		.write_port_out_pel_2(wr_line_buffer_0_2_out_pel.actor),        
		.write_port_out_pel_3(wr_line_buffer_0_3_out_pel.actor),        
		.write_port_out_pel_4(wr_line_buffer_0_4_out_pel.actor),        
		.write_port_out_pel_5(wr_line_buffer_0_5_out_pel.actor),        
		.write_port_out_pel_6(wr_line_buffer_0_6_out_pel.actor),        
		.write_port_out_pel_7(wr_line_buffer_0_7_out_pel.actor)        		
        );

        //line_buffer_1
        line_buffer_8p#(FLUX) line_buffer1
        (
        .clk(clk),
        .rst(rst),        
        .read_port_real_size(rd_line_buffer_1_real_size.actor),
        .read_port_ext_size(rd_line_buffer_1_ext_size.actor),
        .read_port_in_pel_0(rd_line_buffer_1_0_in_pel.actor),            
		.read_port_in_pel_1(rd_line_buffer_1_1_in_pel.actor),            
		.read_port_in_pel_2(rd_line_buffer_1_2_in_pel.actor),            
		.read_port_in_pel_3(rd_line_buffer_1_3_in_pel.actor),            
		.read_port_in_pel_4(rd_line_buffer_1_4_in_pel.actor),            
		.read_port_in_pel_5(rd_line_buffer_1_5_in_pel.actor),            
		.read_port_in_pel_6(rd_line_buffer_1_6_in_pel.actor),            
		.read_port_in_pel_7(rd_line_buffer_1_7_in_pel.actor),
		.write_port_out_pel_0(wr_line_buffer_1_0_out_pel.actor),        		
        .write_port_out_pel_1(wr_line_buffer_1_1_out_pel.actor),        
		.write_port_out_pel_2(wr_line_buffer_1_2_out_pel.actor),        
		.write_port_out_pel_3(wr_line_buffer_1_3_out_pel.actor),        
		.write_port_out_pel_4(wr_line_buffer_1_4_out_pel.actor),        
		.write_port_out_pel_5(wr_line_buffer_1_5_out_pel.actor),        
		.write_port_out_pel_6(wr_line_buffer_1_6_out_pel.actor),        
		.write_port_out_pel_7(wr_line_buffer_1_7_out_pel.actor)        		
        );
               
        //line_buffer_2
        line_buffer_8p#(FLUX) line_buffer2
        (
        .clk(clk),
        .rst(rst),        
        .read_port_real_size(rd_line_buffer_2_real_size.actor),
        .read_port_ext_size(rd_line_buffer_2_ext_size.actor),
        .read_port_in_pel_0(rd_line_buffer_2_0_in_pel.actor),            
		.read_port_in_pel_1(rd_line_buffer_2_1_in_pel.actor),            
		.read_port_in_pel_2(rd_line_buffer_2_2_in_pel.actor),            
		.read_port_in_pel_3(rd_line_buffer_2_3_in_pel.actor),            
		.read_port_in_pel_4(rd_line_buffer_2_4_in_pel.actor),            
		.read_port_in_pel_5(rd_line_buffer_2_5_in_pel.actor),            
		.read_port_in_pel_6(rd_line_buffer_2_6_in_pel.actor),            
		.read_port_in_pel_7(rd_line_buffer_2_7_in_pel.actor),
		.write_port_out_pel_0(wr_line_buffer_2_0_out_pel.actor),        		
        .write_port_out_pel_1(wr_line_buffer_2_1_out_pel.actor),        
		.write_port_out_pel_2(wr_line_buffer_2_2_out_pel.actor),        
		.write_port_out_pel_3(wr_line_buffer_2_3_out_pel.actor),        
		.write_port_out_pel_4(wr_line_buffer_2_4_out_pel.actor),        
		.write_port_out_pel_5(wr_line_buffer_2_5_out_pel.actor),        
		.write_port_out_pel_6(wr_line_buffer_2_6_out_pel.actor),        
		.write_port_out_pel_7(wr_line_buffer_2_7_out_pel.actor)        		
        );

        //line_buffer_3
        line_buffer_8p#(FLUX) line_buffer3
        (
        .clk(clk),
        .rst(rst),        
        .read_port_real_size(rd_line_buffer_3_real_size.actor),
        .read_port_ext_size(rd_line_buffer_3_ext_size.actor),
        .read_port_in_pel_0(rd_line_buffer_3_0_in_pel.actor),            
		.read_port_in_pel_1(rd_line_buffer_3_1_in_pel.actor),            
		.read_port_in_pel_2(rd_line_buffer_3_2_in_pel.actor),            
		.read_port_in_pel_3(rd_line_buffer_3_3_in_pel.actor),            
		.read_port_in_pel_4(rd_line_buffer_3_4_in_pel.actor),            
		.read_port_in_pel_5(rd_line_buffer_3_5_in_pel.actor),            
		.read_port_in_pel_6(rd_line_buffer_3_6_in_pel.actor),            
		.read_port_in_pel_7(rd_line_buffer_3_7_in_pel.actor),
		.write_port_out_pel_0(wr_line_buffer_3_0_out_pel.actor),        		
        .write_port_out_pel_1(wr_line_buffer_3_1_out_pel.actor),        
		.write_port_out_pel_2(wr_line_buffer_3_2_out_pel.actor),        
		.write_port_out_pel_3(wr_line_buffer_3_3_out_pel.actor),        
		.write_port_out_pel_4(wr_line_buffer_3_4_out_pel.actor),        
		.write_port_out_pel_5(wr_line_buffer_3_5_out_pel.actor),        
		.write_port_out_pel_6(wr_line_buffer_3_6_out_pel.actor),        
		.write_port_out_pel_7(wr_line_buffer_3_7_out_pel.actor)        		
        );        
        
        //line_buffer_4
        line_buffer_8p#(FLUX) line_buffer4
        (
        .clk(clk),
        .rst(rst),        
        .read_port_real_size(rd_line_buffer_4_real_size.actor),
        .read_port_ext_size(rd_line_buffer_4_ext_size.actor),
        .read_port_in_pel_0(rd_line_buffer_4_0_in_pel.actor),            
		.read_port_in_pel_1(rd_line_buffer_4_1_in_pel.actor),            
		.read_port_in_pel_2(rd_line_buffer_4_2_in_pel.actor),            
		.read_port_in_pel_3(rd_line_buffer_4_3_in_pel.actor),            
		.read_port_in_pel_4(rd_line_buffer_4_4_in_pel.actor),            
		.read_port_in_pel_5(rd_line_buffer_4_5_in_pel.actor),            
		.read_port_in_pel_6(rd_line_buffer_4_6_in_pel.actor),            
		.read_port_in_pel_7(rd_line_buffer_4_7_in_pel.actor),
		.write_port_out_pel_0(wr_line_buffer_4_0_out_pel.actor),        		
        .write_port_out_pel_1(wr_line_buffer_4_1_out_pel.actor),        
		.write_port_out_pel_2(wr_line_buffer_4_2_out_pel.actor),        
		.write_port_out_pel_3(wr_line_buffer_4_3_out_pel.actor),        
		.write_port_out_pel_4(wr_line_buffer_4_4_out_pel.actor),        
		.write_port_out_pel_5(wr_line_buffer_4_5_out_pel.actor),        
		.write_port_out_pel_6(wr_line_buffer_4_6_out_pel.actor),        
		.write_port_out_pel_7(wr_line_buffer_4_7_out_pel.actor)        		
        );
        
         //line_buffer_5
        line_buffer_8p#(FLUX) line_buffer5
        (
        .clk(clk),
        .rst(rst),        
        .read_port_real_size(rd_line_buffer_5_real_size.actor),
        .read_port_ext_size(rd_line_buffer_5_ext_size.actor),
        .read_port_in_pel_0(rd_line_buffer_5_0_in_pel.actor),            
		.read_port_in_pel_1(rd_line_buffer_5_1_in_pel.actor),            
		.read_port_in_pel_2(rd_line_buffer_5_2_in_pel.actor),            
		.read_port_in_pel_3(rd_line_buffer_5_3_in_pel.actor),            
		.read_port_in_pel_4(rd_line_buffer_5_4_in_pel.actor),            
		.read_port_in_pel_5(rd_line_buffer_5_5_in_pel.actor),            
		.read_port_in_pel_6(rd_line_buffer_5_6_in_pel.actor),            
		.read_port_in_pel_7(rd_line_buffer_5_7_in_pel.actor),
		.write_port_out_pel_0(wr_line_buffer_5_0_out_pel.actor),        		
        .write_port_out_pel_1(wr_line_buffer_5_1_out_pel.actor),        
		.write_port_out_pel_2(wr_line_buffer_5_2_out_pel.actor),        
		.write_port_out_pel_3(wr_line_buffer_5_3_out_pel.actor),        
		.write_port_out_pel_4(wr_line_buffer_5_4_out_pel.actor),        
		.write_port_out_pel_5(wr_line_buffer_5_5_out_pel.actor),        
		.write_port_out_pel_6(wr_line_buffer_5_6_out_pel.actor),        
		.write_port_out_pel_7(wr_line_buffer_5_7_out_pel.actor)        		
        );        
        
        //line_buffer_6
        line_buffer_8p#(FLUX) line_buffer6
        (
        .clk(clk),
        .rst(rst),        
        .read_port_real_size(rd_line_buffer_6_real_size.actor),
        .read_port_ext_size(rd_line_buffer_6_ext_size.actor),
        .read_port_in_pel_0(rd_line_buffer_6_0_in_pel.actor),            
		.read_port_in_pel_1(rd_line_buffer_6_1_in_pel.actor),            
		.read_port_in_pel_2(rd_line_buffer_6_2_in_pel.actor),            
		.read_port_in_pel_3(rd_line_buffer_6_3_in_pel.actor),            
		.read_port_in_pel_4(rd_line_buffer_6_4_in_pel.actor),            
		.read_port_in_pel_5(rd_line_buffer_6_5_in_pel.actor),            
		.read_port_in_pel_6(rd_line_buffer_6_6_in_pel.actor),            
		.read_port_in_pel_7(rd_line_buffer_6_7_in_pel.actor),
		.write_port_out_pel_0(wr_line_buffer_6_0_out_pel.actor),        		
        .write_port_out_pel_1(wr_line_buffer_6_1_out_pel.actor),        
		.write_port_out_pel_2(wr_line_buffer_6_2_out_pel.actor),        
		.write_port_out_pel_3(wr_line_buffer_6_3_out_pel.actor),        
		.write_port_out_pel_4(wr_line_buffer_6_4_out_pel.actor),        
		.write_port_out_pel_5(wr_line_buffer_6_5_out_pel.actor),        
		.write_port_out_pel_6(wr_line_buffer_6_6_out_pel.actor),        
		.write_port_out_pel_7(wr_line_buffer_6_7_out_pel.actor)        		
        ); 
        
    //SHIFT (x8); I: VIOLET - O: FUCSIA

        //shift_0 
        shift #(FLUX) shift_0
        (
        .read_port_in_pel(rd_shift_0_in_pel.actor),    
        .write_port_out_pel(wr_shift_0_out_pel.actor)        
        );

        //shift_1
        shift #(FLUX) shift_1
        (
        .read_port_in_pel(rd_shift_1_in_pel.actor),    
        .write_port_out_pel(wr_shift_1_out_pel.actor)        
        );
        
        //shift_2
        shift #(FLUX) shift_2
        (
        .read_port_in_pel(rd_shift_2_in_pel.actor),    
        .write_port_out_pel(wr_shift_2_out_pel.actor)        
        );		
		
        //shift_3 
        shift #(FLUX) shift_3
        (
        .read_port_in_pel(rd_shift_3_in_pel.actor),    
        .write_port_out_pel(wr_shift_3_out_pel.actor)        
        );
    
        //shift_4
        shift #(FLUX) shift_4
        (
        .read_port_in_pel(rd_shift_4_in_pel.actor),    
        .write_port_out_pel(wr_shift_4_out_pel.actor)        
        );

        //shift_5 
        shift #(FLUX) shift_5
        (
        .read_port_in_pel(rd_shift_5_in_pel.actor),    
        .write_port_out_pel(wr_shift_5_out_pel.actor)        
        );
        
        //shift_6 
        shift #(FLUX) shift_6
        (
        .read_port_in_pel(rd_shift_6_in_pel.actor),    
        .write_port_out_pel(wr_shift_6_out_pel.actor)        
        );		
		
        //shift_7 
        shift #(FLUX) shift_7
        (
        .read_port_in_pel(rd_shift_7_in_pel.actor),    
        .write_port_out_pel(wr_shift_7_out_pel.actor)        
        );		
		
    //CLIP (x8); I: FUCSIA - O: PINK

        //clip_0 
        clip #(FLUX) clip_0
        (
        .read_port_in_pel(rd_clip_0_in_pel.actor),    
        .write_port_out_pel(wr_clip_0_out_pel.actor)        
        );

        //clip_1
        clip #(FLUX) clip_1
        (
        .read_port_in_pel(rd_clip_1_in_pel.actor),    
        .write_port_out_pel(wr_clip_1_out_pel.actor)        
        );

        //clip_2 
        clip #(FLUX) clip_2
        (
        .read_port_in_pel(rd_clip_2_in_pel.actor),    
        .write_port_out_pel(wr_clip_2_out_pel.actor)        
        );
		
		//clip_3
        clip #(FLUX) clip_3
        (
        .read_port_in_pel(rd_clip_3_in_pel.actor),    
        .write_port_out_pel(wr_clip_3_out_pel.actor)        
        );
    
	    //clip_4 
        clip #(FLUX) clip_4
        (
        .read_port_in_pel(rd_clip_4_in_pel.actor),    
        .write_port_out_pel(wr_clip_4_out_pel.actor)        
        );
		
	    //clip_5 
        clip #(FLUX) clip_5
        (
        .read_port_in_pel(rd_clip_5_in_pel.actor),    
        .write_port_out_pel(wr_clip_5_out_pel.actor)        
        );	

	    //clip_6 
        clip #(FLUX) clip_6
        (
        .read_port_in_pel(rd_clip_6_in_pel.actor),    
        .write_port_out_pel(wr_clip_6_out_pel.actor)        
        );
		
	    //clip_7 
        clip #(FLUX) clip_7
        (
        .read_port_in_pel(rd_clip_7_in_pel.actor),    
        .write_port_out_pel(wr_clip_7_out_pel.actor)        
        );
	
    //REMOVE_V (x1); I: PINK / BLUE / BROWN - O: NULL
    
    //REMOVE_v (x8); I: LIME/YELLOW - O: DARK GREY (2�HALF) / RED (2�HALF)

        //remove_v_0
        remove_v #(FLUX) remove_v_0
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_remove_v_0_real_size.actor),        
        .read_port_ext_size(rd_remove_v_0_ext_size.actor),
        .read_port_in_pel(rd_remove_v_0_in_pel.actor),
		.write_port_out_pel(wr_remove_v_0_out_pel.actor)
        );
		
		//remove_v_1
        remove_v #(FLUX) remove_v_1
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_remove_v_1_real_size.actor),
        .read_port_ext_size(rd_remove_v_1_ext_size.actor),
        .read_port_in_pel(rd_remove_v_1_in_pel.actor),
		.write_port_out_pel(wr_remove_v_1_out_pel.actor)
        );
		
		//remove_v_2
        remove_v #(FLUX) remove_v_2
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_remove_v_2_real_size.actor),
        .read_port_ext_size(rd_remove_v_2_ext_size.actor),
        .read_port_in_pel(rd_remove_v_2_in_pel.actor),
		.write_port_out_pel(wr_remove_v_2_out_pel.actor)
        );
		
		//remove_v_3
        remove_v #(FLUX) remove_v_3
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_remove_v_3_real_size.actor),
        .read_port_ext_size(rd_remove_v_3_ext_size.actor),
        .read_port_in_pel(rd_remove_v_3_in_pel.actor),
		.write_port_out_pel(wr_remove_v_3_out_pel.actor)
        );
		
		//remove_v_4
        remove_v #(FLUX) remove_v_4
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_remove_v_4_real_size.actor),
        .read_port_ext_size(rd_remove_v_4_ext_size.actor),
        .read_port_in_pel(rd_remove_v_4_in_pel.actor),
		.write_port_out_pel(wr_remove_v_4_out_pel.actor)
        );
		
		//remove_v_5
        remove_v #(FLUX) remove_v_5
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_remove_v_5_real_size.actor),
        .read_port_ext_size(rd_remove_v_5_ext_size.actor),
        .read_port_in_pel(rd_remove_v_5_in_pel.actor),
		.write_port_out_pel(wr_remove_v_5_out_pel.actor)
        );
		
		//remove_v_6
        remove_v #(FLUX) remove_v_6
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_remove_v_6_real_size.actor),
        .read_port_ext_size(rd_remove_v_6_ext_size.actor),
        .read_port_in_pel(rd_remove_v_6_in_pel.actor),
		.write_port_out_pel(wr_remove_v_6_out_pel.actor)
        );
		
		//remove_v_7
        remove_v #(FLUX) remove_v_7
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_remove_v_7_real_size.actor),
        .read_port_ext_size(rd_remove_v_7_ext_size.actor),
        .read_port_in_pel(rd_remove_v_7_in_pel.actor),
		.write_port_out_pel(wr_remove_v_7_out_pel.actor)
        );
   
      
   //add27 (x56); I: BORDEAUX/GREEN - O: GREEN / YELLOW

	//1� adder tree
    
        //add27_0
        add_27 #(FLUX) add27_0
        (
        .read_port_opA(rd_add_27_0_opA.actor),
        .read_port_opB(rd_add_27_0_opB.actor),    
        .write_port_sum(wr_add_27_0_sum.actor)        
        );
    
        //add27_1 
        add_27 #(FLUX) add27_1 
        (
        .read_port_opA(rd_add_27_1_opA.actor),
        .read_port_opB(rd_add_27_1_opB.actor),    
        .write_port_sum(wr_add_27_1_sum.actor)        
        );
    
        //add27_2
        add_27 #(FLUX) add27_2 
        (
        .read_port_opA(rd_add_27_2_opA.actor),
        .read_port_opB(rd_add_27_2_opB.actor),    
        .write_port_sum(wr_add_27_2_sum.actor)        
        );
    
        //add27_3
        add_27 #(FLUX) add27_3
        (
        .read_port_opA(rd_add_27_3_opA.actor),
        .read_port_opB(rd_add_27_3_opB.actor),    
        .write_port_sum(wr_add_27_3_sum.actor)        
        );
        
        //add27_4 
        add_27 #(FLUX) add27_4 
        (
        .read_port_opA(rd_add_27_4_opA.actor),
        .read_port_opB(rd_add_27_4_opB.actor),    
        .write_port_sum(wr_add_27_4_sum.actor)        
        );
    
        //add27_5 
        add_27 #(FLUX) add27_5 
        (
        .read_port_opA(rd_add_27_5_opA.actor),
        .read_port_opB(rd_add_27_5_opB.actor),    
        .write_port_sum(wr_add_27_5_sum.actor)        
        );
        
        //add27_6
        add_27 #(FLUX) add27_6
        (
        .read_port_opA(rd_add_27_6_opA.actor),
        .read_port_opB(rd_add_27_6_opB.actor),    
        .write_port_sum(wr_add_27_6_sum.actor)        
        );

	//2� adder tree
    
        //add27_7
        add_27 #(FLUX) add27_7
        (
        .read_port_opA(rd_add_27_7_opA.actor),
        .read_port_opB(rd_add_27_7_opB.actor),    
        .write_port_sum(wr_add_27_7_sum.actor)        
        );
    
        //add27_8 
        add_27 #(FLUX) add27_8 
        (
        .read_port_opA(rd_add_27_8_opA.actor),
        .read_port_opB(rd_add_27_8_opB.actor),    
        .write_port_sum(wr_add_27_8_sum.actor)        
        );
    
        //add27_9
        add_27 #(FLUX) add27_9 
        (
        .read_port_opA(rd_add_27_9_opA.actor),
        .read_port_opB(rd_add_27_9_opB.actor),    
        .write_port_sum(wr_add_27_9_sum.actor)        
        );
    
        //add27_10
        add_27 #(FLUX) add27_10
        (
        .read_port_opA(rd_add_27_10_opA.actor),
        .read_port_opB(rd_add_27_10_opB.actor),    
        .write_port_sum(wr_add_27_10_sum.actor)        
        );
        
        //add27_11 
        add_27 #(FLUX) add27_11 
        (
        .read_port_opA(rd_add_27_11_opA.actor),
        .read_port_opB(rd_add_27_11_opB.actor),    
        .write_port_sum(wr_add_27_11_sum.actor)        
        );
    
        //add27_12 
        add_27 #(FLUX) add27_12
        (
        .read_port_opA(rd_add_27_12_opA.actor),
        .read_port_opB(rd_add_27_12_opB.actor),    
        .write_port_sum(wr_add_27_12_sum.actor)        
        );
        
        //add27_13
        add_27 #(FLUX) add27_13
        (
        .read_port_opA(rd_add_27_13_opA.actor),
        .read_port_opB(rd_add_27_13_opB.actor),    
        .write_port_sum(wr_add_27_13_sum.actor)        
        );
		
	//3� adder tree
    
        //add27_14
        add_27 #(FLUX) add27_14
        (
        .read_port_opA(rd_add_27_14_opA.actor),
        .read_port_opB(rd_add_27_14_opB.actor),    
        .write_port_sum(wr_add_27_14_sum.actor)        
        );
    
        //add27_15 
        add_27 #(FLUX) add27_15
        (
        .read_port_opA(rd_add_27_15_opA.actor),
        .read_port_opB(rd_add_27_15_opB.actor),    
        .write_port_sum(wr_add_27_15_sum.actor)        
        );
    
        //add27_16
        add_27 #(FLUX) add27_16
        (
        .read_port_opA(rd_add_27_16_opA.actor),
        .read_port_opB(rd_add_27_16_opB.actor),    
        .write_port_sum(wr_add_27_16_sum.actor)        
        );
    
        //add27_17
        add_27 #(FLUX) add27_17
        (
        .read_port_opA(rd_add_27_17_opA.actor),
        .read_port_opB(rd_add_27_17_opB.actor),    
        .write_port_sum(wr_add_27_17_sum.actor)        
        );
        
        //add27_18 
        add_27 #(FLUX) add27_18
        (
        .read_port_opA(rd_add_27_18_opA.actor),
        .read_port_opB(rd_add_27_18_opB.actor),    
        .write_port_sum(wr_add_27_18_sum.actor)        
        );
    
        //add27_19 
        add_27 #(FLUX) add27_19 
        (
        .read_port_opA(rd_add_27_19_opA.actor),
        .read_port_opB(rd_add_27_19_opB.actor),    
        .write_port_sum(wr_add_27_19_sum.actor)        
        );
        
        //add27_20
        add_27 #(FLUX) add27_20
        (
        .read_port_opA(rd_add_27_20_opA.actor),
        .read_port_opB(rd_add_27_20_opB.actor),    
        .write_port_sum(wr_add_27_20_sum.actor)        
        );		
		
	//4�adder tree
    
        //add27_21
        add_27 #(FLUX) add27_21
        (
        .read_port_opA(rd_add_27_21_opA.actor),
        .read_port_opB(rd_add_27_21_opB.actor),    
        .write_port_sum(wr_add_27_21_sum.actor)        
        );
    
        //add27_22
        add_27 #(FLUX) add27_22
        (
        .read_port_opA(rd_add_27_22_opA.actor),
        .read_port_opB(rd_add_27_22_opB.actor),    
        .write_port_sum(wr_add_27_22_sum.actor)        
        );
    
        //add27_23
        add_27 #(FLUX) add27_23
        (
        .read_port_opA(rd_add_27_23_opA.actor),
        .read_port_opB(rd_add_27_23_opB.actor),    
        .write_port_sum(wr_add_27_23_sum.actor)        
        );
    
        //add27_24
        add_27 #(FLUX) add27_24
        (
        .read_port_opA(rd_add_27_24_opA.actor),
        .read_port_opB(rd_add_27_24_opB.actor),    
        .write_port_sum(wr_add_27_24_sum.actor)        
        );
        
        //add27_25 
        add_27 #(FLUX) add27_25
        (
        .read_port_opA(rd_add_27_25_opA.actor),
        .read_port_opB(rd_add_27_25_opB.actor),    
        .write_port_sum(wr_add_27_25_sum.actor)        
        );
    
        //add27_26 
        add_27 #(FLUX) add27_26
        (
        .read_port_opA(rd_add_27_26_opA.actor),
        .read_port_opB(rd_add_27_26_opB.actor),    
        .write_port_sum(wr_add_27_26_sum.actor)        
        );
        
        //add27_27
        add_27 #(FLUX) add27_27
        (
        .read_port_opA(rd_add_27_27_opA.actor),
        .read_port_opB(rd_add_27_27_opB.actor),    
        .write_port_sum(wr_add_27_27_sum.actor)        
        );

	//5�adder tree
    
        //add27_28
        add_27 #(FLUX) add27_28
        (
        .read_port_opA(rd_add_27_28_opA.actor),
        .read_port_opB(rd_add_27_28_opB.actor),    
        .write_port_sum(wr_add_27_28_sum.actor)        
        );
    
        //add27_29
        add_27 #(FLUX) add27_29
        (
        .read_port_opA(rd_add_27_29_opA.actor),
        .read_port_opB(rd_add_27_29_opB.actor),    
        .write_port_sum(wr_add_27_29_sum.actor)        
        );
    
        //add27_30
        add_27 #(FLUX) add27_30
        (
        .read_port_opA(rd_add_27_30_opA.actor),
        .read_port_opB(rd_add_27_30_opB.actor),    
        .write_port_sum(wr_add_27_30_sum.actor)        
        );
    
        //add27_31
        add_27 #(FLUX) add27_31
        (
        .read_port_opA(rd_add_27_31_opA.actor),
        .read_port_opB(rd_add_27_31_opB.actor),    
        .write_port_sum(wr_add_27_31_sum.actor)        
        );
        
        //add27_32
        add_27 #(FLUX) add27_32
        (
        .read_port_opA(rd_add_27_32_opA.actor),
        .read_port_opB(rd_add_27_32_opB.actor),    
        .write_port_sum(wr_add_27_32_sum.actor)        
        );
    
        //add27_33
        add_27 #(FLUX) add27_33 
        (
        .read_port_opA(rd_add_27_33_opA.actor),
        .read_port_opB(rd_add_27_33_opB.actor),    
        .write_port_sum(wr_add_27_33_sum.actor)        
        );
        
        //add27_34
        add_27 #(FLUX) add27_34
        (
        .read_port_opA(rd_add_27_34_opA.actor),
        .read_port_opB(rd_add_27_34_opB.actor),    
        .write_port_sum(wr_add_27_34_sum.actor)        
        );

	//6�adder tree
    
        //add27_35
        add_27 #(FLUX) add27_35
        (
        .read_port_opA(rd_add_27_35_opA.actor),
        .read_port_opB(rd_add_27_35_opB.actor),    
        .write_port_sum(wr_add_27_35_sum.actor)        
        );
    
        //add27_36 
        add_27 #(FLUX) add27_36 
        (
        .read_port_opA(rd_add_27_36_opA.actor),
        .read_port_opB(rd_add_27_36_opB.actor),    
        .write_port_sum(wr_add_27_36_sum.actor)        
        );
    
        //add27_37
        add_27 #(FLUX) add27_37
        (
        .read_port_opA(rd_add_27_37_opA.actor),
        .read_port_opB(rd_add_27_37_opB.actor),    
        .write_port_sum(wr_add_27_37_sum.actor)        
        );
    
        //add27_38
        add_27 #(FLUX) add27_38
        (
        .read_port_opA(rd_add_27_38_opA.actor),
        .read_port_opB(rd_add_27_38_opB.actor),    
        .write_port_sum(wr_add_27_38_sum.actor)        
        );
        
        //add27_39 
        add_27 #(FLUX) add27_39
        (
        .read_port_opA(rd_add_27_39_opA.actor),
        .read_port_opB(rd_add_27_39_opB.actor),    
        .write_port_sum(wr_add_27_39_sum.actor)        
        );
    
        //add27_40 
        add_27 #(FLUX) add27_40
        (
        .read_port_opA(rd_add_27_40_opA.actor),
        .read_port_opB(rd_add_27_40_opB.actor),    
        .write_port_sum(wr_add_27_40_sum.actor)        
        );
        
        //add27_41
        add_27 #(FLUX) add27_41
        (
        .read_port_opA(rd_add_27_41_opA.actor),
        .read_port_opB(rd_add_27_41_opB.actor),    
        .write_port_sum(wr_add_27_41_sum.actor)        
        );
        
	//7�adder tree
    
        //add27_42
        add_27 #(FLUX) add27_42
        (
        .read_port_opA(rd_add_27_42_opA.actor),
        .read_port_opB(rd_add_27_42_opB.actor),    
        .write_port_sum(wr_add_27_42_sum.actor)        
        );
    
        //add27_43 
        add_27 #(FLUX) add27_43 
        (
        .read_port_opA(rd_add_27_43_opA.actor),
        .read_port_opB(rd_add_27_43_opB.actor),    
        .write_port_sum(wr_add_27_43_sum.actor)        
        );
    
        //add27_44
        add_27 #(FLUX) add27_44
        (
        .read_port_opA(rd_add_27_44_opA.actor),
        .read_port_opB(rd_add_27_44_opB.actor),    
        .write_port_sum(wr_add_27_44_sum.actor)        
        );
    
        //add27_45
        add_27 #(FLUX) add27_45
        (
        .read_port_opA(rd_add_27_45_opA.actor),
        .read_port_opB(rd_add_27_45_opB.actor),    
        .write_port_sum(wr_add_27_45_sum.actor)        
        );
        
        //add27_46 
        add_27 #(FLUX) add27_46 
        (
        .read_port_opA(rd_add_27_46_opA.actor),
        .read_port_opB(rd_add_27_46_opB.actor),    
        .write_port_sum(wr_add_27_46_sum.actor)        
        );
    
        //add27_47 
        add_27 #(FLUX) add27_47 
        (
        .read_port_opA(rd_add_27_47_opA.actor),
        .read_port_opB(rd_add_27_47_opB.actor),    
        .write_port_sum(wr_add_27_47_sum.actor)        
        );
        
        //add27_48
        add_27 #(FLUX) add27_48
        (
        .read_port_opA(rd_add_27_48_opA.actor),
        .read_port_opB(rd_add_27_48_opB.actor),    
        .write_port_sum(wr_add_27_48_sum.actor)        
        );

	//8� adder tree
    
        //add27_49
        add_27 #(FLUX) add27_49
        (
        .read_port_opA(rd_add_27_49_opA.actor),
        .read_port_opB(rd_add_27_49_opB.actor),    
        .write_port_sum(wr_add_27_49_sum.actor)        
        );
    
        //add27_50
        add_27 #(FLUX) add27_50 
        (
        .read_port_opA(rd_add_27_50_opA.actor),
        .read_port_opB(rd_add_27_50_opB.actor),    
        .write_port_sum(wr_add_27_50_sum.actor)        
        );
    
        //add27_51
        add_27 #(FLUX) add27_51
        (
        .read_port_opA(rd_add_27_51_opA.actor),
        .read_port_opB(rd_add_27_51_opB.actor),    
        .write_port_sum(wr_add_27_51_sum.actor)        
        );
    
        //add27_52
        add_27 #(FLUX) add27_52
        (
        .read_port_opA(rd_add_27_52_opA.actor),
        .read_port_opB(rd_add_27_52_opB.actor),    
        .write_port_sum(wr_add_27_52_sum.actor)        
        );
        
        //add27_53 
        add_27 #(FLUX) add27_53 
        (
        .read_port_opA(rd_add_27_53_opA.actor),
        .read_port_opB(rd_add_27_53_opB.actor),    
        .write_port_sum(wr_add_27_53_sum.actor)        
        );
    
        //add27_54 
        add_27 #(FLUX) add27_54 
        (
        .read_port_opA(rd_add_27_54_opA.actor),
        .read_port_opB(rd_add_27_54_opB.actor),    
        .write_port_sum(wr_add_27_54_sum.actor)        
        );
        
        //add27_55
        add_27 #(FLUX) add27_55
        (
        .read_port_opA(rd_add_27_55_opA.actor),
        .read_port_opB(rd_add_27_55_opB.actor),    
        .write_port_sum(wr_add_27_55_sum.actor)        
        );
		
    //mul18 (x64); I: DARK YELLOW/RED/BEIGE - O: BORDEAUX / GREEN
    
	//1� colonna
	
        //mul18_0
        mul_18 #(FLUX) mul18_0
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_0_real_size.actor),
        .read_port_ext_size(rd_mul_18_0_ext_size.actor),
        .read_port_opA(rd_mul_18_0_opA.actor),
        .read_port_opB(rd_mul_18_0_opB.actor),        
        .write_port_prod(wr_mul_18_0_prod.actor)        
        );
    
        //mul18_1
        mul_18 #(FLUX) mul18_1
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_1_real_size.actor),
        .read_port_ext_size(rd_mul_18_1_ext_size.actor),
        .read_port_opA(rd_mul_18_1_opA.actor),
        .read_port_opB(rd_mul_18_1_opB.actor),        
        .write_port_prod(wr_mul_18_1_prod.actor)        
        );
    
        //mul18_2
        mul_18 #(FLUX) mul18_2
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_2_real_size.actor),
        .read_port_ext_size(rd_mul_18_2_ext_size.actor),
        .read_port_opA(rd_mul_18_2_opA.actor),
        .read_port_opB(rd_mul_18_2_opB.actor),        
        .write_port_prod(wr_mul_18_2_prod.actor)        
        );
    
        //mul18_3
        mul_18 #(FLUX) mul18_3
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_3_real_size.actor),
        .read_port_ext_size(rd_mul_18_3_ext_size.actor),
        .read_port_opA(rd_mul_18_3_opA.actor),
        .read_port_opB(rd_mul_18_3_opB.actor),        
        .write_port_prod(wr_mul_18_3_prod.actor)        
        );
    
        //mul18_4
        mul_18 #(FLUX) mul18_4
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_4_real_size.actor),
        .read_port_ext_size(rd_mul_18_4_ext_size.actor),
        .read_port_opA(rd_mul_18_4_opA.actor),
        .read_port_opB(rd_mul_18_4_opB.actor),        
        .write_port_prod(wr_mul_18_4_prod.actor)        
        );
    
        //mul18_5
        mul_18 #(FLUX) mul18_5
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_5_real_size.actor),
        .read_port_ext_size(rd_mul_18_5_ext_size.actor),
        .read_port_opA(rd_mul_18_5_opA.actor),
        .read_port_opB(rd_mul_18_5_opB.actor),        
        .write_port_prod(wr_mul_18_5_prod.actor)        
        );
    
        //mul18_6
        mul_18 #(FLUX) mul18_6
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_6_real_size.actor),
        .read_port_ext_size(rd_mul_18_6_ext_size.actor),
        .read_port_opA(rd_mul_18_6_opA.actor),
        .read_port_opB(rd_mul_18_6_opB.actor),        
        .write_port_prod(wr_mul_18_6_prod.actor)        
        );
    
        //mul18_7
        mul_18 #(FLUX) mul18_7
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_7_real_size.actor),
        .read_port_ext_size(rd_mul_18_7_ext_size.actor),
        .read_port_opA(rd_mul_18_7_opA.actor),
        .read_port_opB(rd_mul_18_7_opB.actor),        
        .write_port_prod(wr_mul_18_7_prod.actor)        
        );
    
	//2� colonna

        //mul18_8
        mul_18 #(FLUX) mul18_8
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_8_real_size.actor),
        .read_port_ext_size(rd_mul_18_8_ext_size.actor),
        .read_port_opA(rd_mul_18_8_opA.actor),
        .read_port_opB(rd_mul_18_8_opB.actor),        
        .write_port_prod(wr_mul_18_8_prod.actor)        
        );

        //mul18_9
        mul_18 #(FLUX) mul18_9
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_9_real_size.actor),
        .read_port_ext_size(rd_mul_18_9_ext_size.actor),
        .read_port_opA(rd_mul_18_9_opA.actor),
        .read_port_opB(rd_mul_18_9_opB.actor),        
        .write_port_prod(wr_mul_18_9_prod.actor)        
        );
    
        //mul18_10
        mul_18 #(FLUX) mul18_10
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_10_real_size.actor),
        .read_port_ext_size(rd_mul_18_10_ext_size.actor),
        .read_port_opA(rd_mul_18_10_opA.actor),
        .read_port_opB(rd_mul_18_10_opB.actor),        
        .write_port_prod(wr_mul_18_10_prod.actor)        
        );
    
        //mul18_11
        mul_18 #(FLUX) mul18_11
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_11_real_size.actor),
        .read_port_ext_size(rd_mul_18_11_ext_size.actor),
        .read_port_opA(rd_mul_18_11_opA.actor),
        .read_port_opB(rd_mul_18_11_opB.actor),        
        .write_port_prod(wr_mul_18_11_prod.actor)        
        );
    
        //mul18_12
        mul_18 #(FLUX) mul18_12
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_12_real_size.actor),
        .read_port_ext_size(rd_mul_18_12_ext_size.actor),
        .read_port_opA(rd_mul_18_12_opA.actor),
        .read_port_opB(rd_mul_18_12_opB.actor),        
        .write_port_prod(wr_mul_18_12_prod.actor)        
        );
    
        //mul18_13
        mul_18 #(FLUX) mul18_13
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_13_real_size.actor),
        .read_port_ext_size(rd_mul_18_13_ext_size.actor),
        .read_port_opA(rd_mul_18_13_opA.actor),
        .read_port_opB(rd_mul_18_13_opB.actor),        
        .write_port_prod(wr_mul_18_13_prod.actor)        
        );
    
        //mul18_14
        mul_18 #(FLUX) mul18_14
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_14_real_size.actor),
        .read_port_ext_size(rd_mul_18_14_ext_size.actor),
        .read_port_opA(rd_mul_18_14_opA.actor),
        .read_port_opB(rd_mul_18_14_opB.actor),        
        .write_port_prod(wr_mul_18_14_prod.actor)        
        );
        
        //mul18_15
        mul_18 #(FLUX) mul18_15
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_15_real_size.actor),
        .read_port_ext_size(rd_mul_18_15_ext_size.actor),
        .read_port_opA(rd_mul_18_15_opA.actor),
        .read_port_opB(rd_mul_18_15_opB.actor),        
        .write_port_prod(wr_mul_18_15_prod.actor)        
        );
		
	//3�colonna

        //mul18_16
        mul_18 #(FLUX) mul18_16
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_16_real_size.actor),
        .read_port_ext_size(rd_mul_18_16_ext_size.actor),
        .read_port_opA(rd_mul_18_16_opA.actor),
        .read_port_opB(rd_mul_18_16_opB.actor),        
        .write_port_prod(wr_mul_18_16_prod.actor)        
        );
    
        //mul18_17
        mul_18 #(FLUX) mul18_17
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_17_real_size.actor),
        .read_port_ext_size(rd_mul_18_17_ext_size.actor),
        .read_port_opA(rd_mul_18_17_opA.actor),
        .read_port_opB(rd_mul_18_17_opB.actor),        
        .write_port_prod(wr_mul_18_17_prod.actor)        
        );
    
        //mul18_18
        mul_18 #(FLUX) mul18_18
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_18_real_size.actor),
        .read_port_ext_size(rd_mul_18_18_ext_size.actor),
        .read_port_opA(rd_mul_18_18_opA.actor),
        .read_port_opB(rd_mul_18_18_opB.actor),        
        .write_port_prod(wr_mul_18_18_prod.actor)        
        );
    
        //mul18_19
        mul_18 #(FLUX) mul18_19
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_19_real_size.actor),
        .read_port_ext_size(rd_mul_18_19_ext_size.actor),
        .read_port_opA(rd_mul_18_19_opA.actor),
        .read_port_opB(rd_mul_18_19_opB.actor),        
        .write_port_prod(wr_mul_18_19_prod.actor)        
        );
    
        //mul18_20
        mul_18 #(FLUX) mul18_20
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_20_real_size.actor),
        .read_port_ext_size(rd_mul_18_20_ext_size.actor),
        .read_port_opA(rd_mul_18_20_opA.actor),
        .read_port_opB(rd_mul_18_20_opB.actor),        
        .write_port_prod(wr_mul_18_20_prod.actor)        
        );
    
        //mul18_21
        mul_18 #(FLUX) mul18_21
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_21_real_size.actor),
        .read_port_ext_size(rd_mul_18_21_ext_size.actor),
        .read_port_opA(rd_mul_18_21_opA.actor),
        .read_port_opB(rd_mul_18_21_opB.actor),        
        .write_port_prod(wr_mul_18_21_prod.actor)        
        );
    
        //mul18_22
        mul_18 #(FLUX) mul18_22
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_22_real_size.actor),
        .read_port_ext_size(rd_mul_18_22_ext_size.actor),
        .read_port_opA(rd_mul_18_22_opA.actor),
        .read_port_opB(rd_mul_18_22_opB.actor),        
        .write_port_prod(wr_mul_18_22_prod.actor)        
        );
    
        //mul18_23
        mul_18 #(FLUX) mul18_23
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_23_real_size.actor),
        .read_port_ext_size(rd_mul_18_23_ext_size.actor),
        .read_port_opA(rd_mul_18_23_opA.actor),
        .read_port_opB(rd_mul_18_23_opB.actor),        
        .write_port_prod(wr_mul_18_23_prod.actor)        
        );
		
	//4�colonna

        //mul18_24
        mul_18 #(FLUX) mul18_24
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_24_real_size.actor),
        .read_port_ext_size(rd_mul_18_24_ext_size.actor),
        .read_port_opA(rd_mul_18_24_opA.actor),
        .read_port_opB(rd_mul_18_24_opB.actor),        
        .write_port_prod(wr_mul_18_24_prod.actor)        
        );
    
        //mul18_25
        mul_18 #(FLUX) mul18_25
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_25_real_size.actor),
        .read_port_ext_size(rd_mul_18_25_ext_size.actor),
        .read_port_opA(rd_mul_18_25_opA.actor),
        .read_port_opB(rd_mul_18_25_opB.actor),        
        .write_port_prod(wr_mul_18_25_prod.actor)        
        );
    
        //mul18_26
        mul_18 #(FLUX) mul18_26
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_26_real_size.actor),
        .read_port_ext_size(rd_mul_18_26_ext_size.actor),
        .read_port_opA(rd_mul_18_26_opA.actor),
        .read_port_opB(rd_mul_18_26_opB.actor),        
        .write_port_prod(wr_mul_18_26_prod.actor)        
        );
    
        //mul18_27
        mul_18 #(FLUX) mul18_27
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_27_real_size.actor),
        .read_port_ext_size(rd_mul_18_27_ext_size.actor),
        .read_port_opA(rd_mul_18_27_opA.actor),
        .read_port_opB(rd_mul_18_27_opB.actor),        
        .write_port_prod(wr_mul_18_27_prod.actor)        
        );
    
        //mul18_28
        mul_18 #(FLUX) mul18_28
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_28_real_size.actor),
        .read_port_ext_size(rd_mul_18_28_ext_size.actor),
        .read_port_opA(rd_mul_18_28_opA.actor),
        .read_port_opB(rd_mul_18_28_opB.actor),        
        .write_port_prod(wr_mul_18_28_prod.actor)        
        );
    
        //mul18_29
        mul_18 #(FLUX) mul18_29
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_29_real_size.actor),
        .read_port_ext_size(rd_mul_18_29_ext_size.actor),
        .read_port_opA(rd_mul_18_29_opA.actor),
        .read_port_opB(rd_mul_18_29_opB.actor),        
        .write_port_prod(wr_mul_18_29_prod.actor)        
        );
    
        //mul18_30
        mul_18 #(FLUX) mul18_30
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_30_real_size.actor),
        .read_port_ext_size(rd_mul_18_30_ext_size.actor),
        .read_port_opA(rd_mul_18_30_opA.actor),
        .read_port_opB(rd_mul_18_30_opB.actor),        
        .write_port_prod(wr_mul_18_30_prod.actor)        
        );
    
        //mul18_31
        mul_18 #(FLUX) mul18_31
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_31_real_size.actor),
        .read_port_ext_size(rd_mul_18_31_ext_size.actor),
        .read_port_opA(rd_mul_18_31_opA.actor),
        .read_port_opB(rd_mul_18_31_opB.actor),        
        .write_port_prod(wr_mul_18_31_prod.actor)        
        );
		
	//5�colonna

        //mul18_32
        mul_18 #(FLUX) mul18_32
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_32_real_size.actor),
        .read_port_ext_size(rd_mul_18_32_ext_size.actor),
        .read_port_opA(rd_mul_18_32_opA.actor),
        .read_port_opB(rd_mul_18_32_opB.actor),        
        .write_port_prod(wr_mul_18_32_prod.actor)        
        );
    
        //mul18_33
        mul_18 #(FLUX) mul18_33
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_33_real_size.actor),
        .read_port_ext_size(rd_mul_18_33_ext_size.actor),
        .read_port_opA(rd_mul_18_33_opA.actor),
        .read_port_opB(rd_mul_18_33_opB.actor),        
        .write_port_prod(wr_mul_18_33_prod.actor)        
        );
    
        //mul18_34
        mul_18 #(FLUX) mul18_34
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_34_real_size.actor),
        .read_port_ext_size(rd_mul_18_34_ext_size.actor),
        .read_port_opA(rd_mul_18_34_opA.actor),
        .read_port_opB(rd_mul_18_34_opB.actor),        
        .write_port_prod(wr_mul_18_34_prod.actor)        
        );
    
        //mul18_35
        mul_18 #(FLUX) mul18_35
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_35_real_size.actor),
        .read_port_ext_size(rd_mul_18_35_ext_size.actor),
        .read_port_opA(rd_mul_18_35_opA.actor),
        .read_port_opB(rd_mul_18_35_opB.actor),        
        .write_port_prod(wr_mul_18_35_prod.actor)        
        );
    
        //mul18_36
        mul_18 #(FLUX) mul18_36
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_36_real_size.actor),
        .read_port_ext_size(rd_mul_18_36_ext_size.actor),
        .read_port_opA(rd_mul_18_36_opA.actor),
        .read_port_opB(rd_mul_18_36_opB.actor),        
        .write_port_prod(wr_mul_18_36_prod.actor)        
        );
    
        //mul18_37
        mul_18 #(FLUX) mul18_37
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_37_real_size.actor),
        .read_port_ext_size(rd_mul_18_37_ext_size.actor),
        .read_port_opA(rd_mul_18_37_opA.actor),
        .read_port_opB(rd_mul_18_37_opB.actor),        
        .write_port_prod(wr_mul_18_37_prod.actor)        
        );
    
        //mul18_38
        mul_18 #(FLUX) mul18_38
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_38_real_size.actor),
        .read_port_ext_size(rd_mul_18_38_ext_size.actor),
        .read_port_opA(rd_mul_18_38_opA.actor),
        .read_port_opB(rd_mul_18_38_opB.actor),        
        .write_port_prod(wr_mul_18_38_prod.actor)        
        );
    
        //mul18_39
        mul_18 #(FLUX) mul18_39
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_39_real_size.actor),
        .read_port_ext_size(rd_mul_18_39_ext_size.actor),
        .read_port_opA(rd_mul_18_39_opA.actor),
        .read_port_opB(rd_mul_18_39_opB.actor),        
        .write_port_prod(wr_mul_18_39_prod.actor)        
        );
		
	//6�colonna

        //mul18_40
        mul_18 #(FLUX) mul18_40
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_40_real_size.actor),
        .read_port_ext_size(rd_mul_18_40_ext_size.actor),
        .read_port_opA(rd_mul_18_40_opA.actor),
        .read_port_opB(rd_mul_18_40_opB.actor),        
        .write_port_prod(wr_mul_18_40_prod.actor)        
        );
    
        //mul18_41
        mul_18 #(FLUX) mul18_41
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_41_real_size.actor),
        .read_port_ext_size(rd_mul_18_41_ext_size.actor),
        .read_port_opA(rd_mul_18_41_opA.actor),
        .read_port_opB(rd_mul_18_41_opB.actor),        
        .write_port_prod(wr_mul_18_41_prod.actor)        
        );
    
        //mul18_42
        mul_18 #(FLUX) mul18_42
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_42_real_size.actor),
        .read_port_ext_size(rd_mul_18_42_ext_size.actor),
        .read_port_opA(rd_mul_18_42_opA.actor),
        .read_port_opB(rd_mul_18_42_opB.actor),        
        .write_port_prod(wr_mul_18_42_prod.actor)        
        );
    
        //mul18_43
        mul_18 #(FLUX) mul18_43
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_43_real_size.actor),
        .read_port_ext_size(rd_mul_18_43_ext_size.actor),
        .read_port_opA(rd_mul_18_43_opA.actor),
        .read_port_opB(rd_mul_18_43_opB.actor),        
        .write_port_prod(wr_mul_18_43_prod.actor)        
        );
    
        //mul18_44
        mul_18 #(FLUX) mul18_44
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_44_real_size.actor),
        .read_port_ext_size(rd_mul_18_44_ext_size.actor),
        .read_port_opA(rd_mul_18_44_opA.actor),
        .read_port_opB(rd_mul_18_44_opB.actor),        
        .write_port_prod(wr_mul_18_44_prod.actor)        
        );
    
        //mul18_45
        mul_18 #(FLUX) mul18_45
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_45_real_size.actor),
        .read_port_ext_size(rd_mul_18_45_ext_size.actor),
        .read_port_opA(rd_mul_18_45_opA.actor),
        .read_port_opB(rd_mul_18_45_opB.actor),        
        .write_port_prod(wr_mul_18_45_prod.actor)        
        );
    
        //mul18_46
        mul_18 #(FLUX) mul18_46
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_46_real_size.actor),
        .read_port_ext_size(rd_mul_18_46_ext_size.actor),
        .read_port_opA(rd_mul_18_46_opA.actor),
        .read_port_opB(rd_mul_18_46_opB.actor),        
        .write_port_prod(wr_mul_18_46_prod.actor)        
        );
    
        //mul18_47
        mul_18 #(FLUX) mul18_47
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_47_real_size.actor),
        .read_port_ext_size(rd_mul_18_47_ext_size.actor),
        .read_port_opA(rd_mul_18_47_opA.actor),
        .read_port_opB(rd_mul_18_47_opB.actor),        
        .write_port_prod(wr_mul_18_47_prod.actor)        
        );
		
	//7�colonna

        //mul18_48
        mul_18 #(FLUX) mul18_48
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_48_real_size.actor),
        .read_port_ext_size(rd_mul_18_48_ext_size.actor),
        .read_port_opA(rd_mul_18_48_opA.actor),
        .read_port_opB(rd_mul_18_48_opB.actor),        
        .write_port_prod(wr_mul_18_48_prod.actor)        
        );
    
        //mul18_49
        mul_18 #(FLUX) mul18_49
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_49_real_size.actor),
        .read_port_ext_size(rd_mul_18_49_ext_size.actor),
        .read_port_opA(rd_mul_18_49_opA.actor),
        .read_port_opB(rd_mul_18_49_opB.actor),        
        .write_port_prod(wr_mul_18_49_prod.actor)        
        );
    
        //mul18_50
        mul_18 #(FLUX) mul18_50
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_50_real_size.actor),
        .read_port_ext_size(rd_mul_18_50_ext_size.actor),
        .read_port_opA(rd_mul_18_50_opA.actor),
        .read_port_opB(rd_mul_18_50_opB.actor),        
        .write_port_prod(wr_mul_18_50_prod.actor)        
        );
    
        //mul18_51
        mul_18 #(FLUX) mul18_51
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_51_real_size.actor),
        .read_port_ext_size(rd_mul_18_51_ext_size.actor),
        .read_port_opA(rd_mul_18_51_opA.actor),
        .read_port_opB(rd_mul_18_51_opB.actor),        
        .write_port_prod(wr_mul_18_51_prod.actor)        
        );
    
        //mul18_52
        mul_18 #(FLUX) mul18_52
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_52_real_size.actor),
        .read_port_ext_size(rd_mul_18_52_ext_size.actor),
        .read_port_opA(rd_mul_18_52_opA.actor),
        .read_port_opB(rd_mul_18_52_opB.actor),        
        .write_port_prod(wr_mul_18_52_prod.actor)        
        );
    
        //mul18_53
        mul_18 #(FLUX) mul18_53
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_53_real_size.actor),
        .read_port_ext_size(rd_mul_18_53_ext_size.actor),
        .read_port_opA(rd_mul_18_53_opA.actor),
        .read_port_opB(rd_mul_18_53_opB.actor),        
        .write_port_prod(wr_mul_18_53_prod.actor)        
        );
    
        //mul18_54
        mul_18 #(FLUX) mul18_54
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_54_real_size.actor),
        .read_port_ext_size(rd_mul_18_54_ext_size.actor),
        .read_port_opA(rd_mul_18_54_opA.actor),
        .read_port_opB(rd_mul_18_54_opB.actor),        
        .write_port_prod(wr_mul_18_54_prod.actor)        
        );
    
        //mul18_55
        mul_18 #(FLUX) mul18_55
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_55_real_size.actor),
        .read_port_ext_size(rd_mul_18_55_ext_size.actor),
        .read_port_opA(rd_mul_18_55_opA.actor),
        .read_port_opB(rd_mul_18_55_opB.actor),        
        .write_port_prod(wr_mul_18_55_prod.actor)        
        );
		
	//8�colonna

        //mul18_56
        mul_18 #(FLUX) mul18_56
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_56_real_size.actor),
        .read_port_ext_size(rd_mul_18_56_ext_size.actor),
        .read_port_opA(rd_mul_18_56_opA.actor),
        .read_port_opB(rd_mul_18_56_opB.actor),        
        .write_port_prod(wr_mul_18_56_prod.actor)        
        );
    
        //mul18_57
        mul_18 #(FLUX) mul18_57
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_57_real_size.actor),
        .read_port_ext_size(rd_mul_18_57_ext_size.actor),
        .read_port_opA(rd_mul_18_57_opA.actor),
        .read_port_opB(rd_mul_18_57_opB.actor),        
        .write_port_prod(wr_mul_18_57_prod.actor)        
        );
    
        //mul18_58
        mul_18 #(FLUX) mul18_58
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_58_real_size.actor),
        .read_port_ext_size(rd_mul_18_58_ext_size.actor),
        .read_port_opA(rd_mul_18_58_opA.actor),
        .read_port_opB(rd_mul_18_58_opB.actor),        
        .write_port_prod(wr_mul_18_58_prod.actor)        
        );
    
        //mul18_59
        mul_18 #(FLUX) mul18_59
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_59_real_size.actor),
        .read_port_ext_size(rd_mul_18_59_ext_size.actor),
        .read_port_opA(rd_mul_18_59_opA.actor),
        .read_port_opB(rd_mul_18_59_opB.actor),        
        .write_port_prod(wr_mul_18_59_prod.actor)        
        );
    
        //mul18_60
        mul_18 #(FLUX) mul18_60
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_60_real_size.actor),
        .read_port_ext_size(rd_mul_18_60_ext_size.actor),
        .read_port_opA(rd_mul_18_60_opA.actor),
        .read_port_opB(rd_mul_18_60_opB.actor),        
        .write_port_prod(wr_mul_18_60_prod.actor)        
        );
    
        //mul18_61
        mul_18 #(FLUX) mul18_61
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_61_real_size.actor),
        .read_port_ext_size(rd_mul_18_61_ext_size.actor),
        .read_port_opA(rd_mul_18_61_opA.actor),
        .read_port_opB(rd_mul_18_61_opB.actor),        
        .write_port_prod(wr_mul_18_61_prod.actor)        
        );
    
        //mul18_62
        mul_18 #(FLUX) mul18_62
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_62_real_size.actor),  
        .read_port_ext_size(rd_mul_18_62_ext_size.actor),
        .read_port_opA(rd_mul_18_62_opA.actor),
        .read_port_opB(rd_mul_18_62_opB.actor),        
        .write_port_prod(wr_mul_18_62_prod.actor)        
        );
    
        //mul18_63
        mul_18 #(FLUX) mul18_63
        (
        .clk(clk),
        .rst(rst),
        .read_port_real_size(rd_mul_18_63_real_size.actor),
        .read_port_ext_size(rd_mul_18_63_ext_size.actor),
        .read_port_opA(rd_mul_18_63_opA.actor),
        .read_port_opB(rd_mul_18_63_opB.actor),        
        .write_port_prod(wr_mul_18_63_prod.actor)        
        );			



//FINE MODULI SECONDA PARTE




//ASSIGN REMOVE_V <-> SEGNALI DI USCITA
     
        assign wr_remove_v_0_out_pel.full=write_port_out_port_0.full;
        assign write_port_out_port_0.write = wr_remove_v_0_out_pel.write;
        assign write_port_out_port_0.din = wr_remove_v_0_out_pel.din;
		
        assign wr_remove_v_1_out_pel.full=write_port_out_port_1.full;
        assign write_port_out_port_1.write = wr_remove_v_1_out_pel.write;
        assign write_port_out_port_1.din = wr_remove_v_1_out_pel.din;		

        assign wr_remove_v_2_out_pel.full=write_port_out_port_2.full;
        assign write_port_out_port_2.write = wr_remove_v_2_out_pel.write;
        assign write_port_out_port_2.din = wr_remove_v_2_out_pel.din;

        assign wr_remove_v_3_out_pel.full=write_port_out_port_3.full;
        assign write_port_out_port_3.write = wr_remove_v_3_out_pel.write;
        assign write_port_out_port_3.din = wr_remove_v_3_out_pel.din;

        assign wr_remove_v_4_out_pel.full=write_port_out_port_4.full;
        assign write_port_out_port_4.write = wr_remove_v_4_out_pel.write;
        assign write_port_out_port_4.din = wr_remove_v_4_out_pel.din;

        assign wr_remove_v_5_out_pel.full=write_port_out_port_5.full;
        assign write_port_out_port_5.write = wr_remove_v_5_out_pel.write;
        assign write_port_out_port_5.din = wr_remove_v_5_out_pel.din;
		
        assign wr_remove_v_6_out_pel.full=write_port_out_port_6.full;
        assign write_port_out_port_6.write = wr_remove_v_6_out_pel.write;
        assign write_port_out_port_6.din = wr_remove_v_6_out_pel.din;		

        assign wr_remove_v_7_out_pel.full=write_port_out_port_7.full;
        assign write_port_out_port_7.write = wr_remove_v_7_out_pel.write;
        assign write_port_out_port_7.din = wr_remove_v_7_out_pel.din;


endmodule